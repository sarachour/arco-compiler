
*constant value 1
Icst4		13	0	DC	1.
*
*@output ES
Vout_ES_3		13	0	DC	1.
*
*@input ES_0
Vin_ES_0_2		13	0	DC	1.
*
*constant value 0.11
Vcst1		12	0	DC	0.11
*
*constant value 0.15
Vcst0		11	0	DC	0.15
*
*
*
* === Connectivity Schem ==== 
XinputI_1		13	10	iin
XoutputV_53		13	0	vout
Xmm_1		3	7	10	10	8	0	0	7	mm
XinputV_1		13	7	vin
XinputV_19		11	3	vin
XinputV_1		13	7	vin
