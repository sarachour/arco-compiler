EXAMPLE PSpice
*
* ## Dependencies
*
.INCLUDE math/basic.subckt
*
* ## Structure
*
VIN1 1 0 DC 2
VIN2 2 0 DC 3

x1 1 2 3 vadd
x2 2 3 4 vmul
*x3 4 1 5 vdiv

*
* ## Analysis and Plotting
*
.OP
.DC
.TF
.DISPLAY
.PLOT x2 V(1)
.END
