
*constant value 0.0008
Vcst55		72	0	DC	0.0008
*
*@input C_0
Vin_C_0_52		72	0	DC	1.
*
*@input DAp_0
Vin_DAp_0_50		71	0	DC	1.
*
*constant value 250
Vcst49		71	0	DC	250.
*
*@input A_0
Vin_A_0_48		70	0	DC	1.
*
*constant value 1
Icst47		70	0	DC	1.
*
*constant value 125
Vcst44		70	0	DC	125.
*
*@input MR_0
Vin_MR_0_43		70	0	DC	1.
*
*constant value 1
Vcst42		69	0	DC	1.
*
*constant value 0.004
Vcst41		69	0	DC	0.004
*
*@input MA_0
Vin_MA_0_40		68	0	DC	1.
*
*constant value 0.2
Icst39		68	0	DC	0.2
*
*@input R_0
Vin_R_0_36		67	0	DC	1.
*
*constant value 0.0204081632653
Icst33		67	0	DC	0.0204081632653
*
*constant value 50
Vcst32		66	0	DC	50.
*
*@input DA_0
Vin_DA_0_31		66	0	DC	1.
*
*constant value 100
Icst30		66	0	DC	100.
*
*constant value -1
Vcst27		66	0	DC	-1.
*
*constant value 0.5
Icst26		66	0	DC	0.5
*
*constant value 500
Icst25		66	0	DC	500.
*
*constant value 100
Vcst24		65	0	DC	100.
*
*@input DR_0
Vin_DR_0_23		64	0	DC	1.
*
*constant value -10
Icst22		64	0	DC	-10.
*
*@input DRp_0
Vin_DRp_0_20		64	0	DC	1.
*
*constant value 0
Icst19		64	0	DC	0.
*
*constant value 10
Icst14		64	0	DC	10.
*
*constant value 0
Vcst12		64	0	DC	0.
*
*constant value 1250
Vcst7		63	0	DC	1250.
*
*constant value 10
Vcst5		62	0	DC	10.
*
*constant value -2500
Vcst4		61	0	DC	-2500.
*
*constant value 0.010101010101
Icst2		60	0	DC	0.010101010101
*
*
*
* === Connectivity Schem ==== 
Xvgain_33		60	60	0	60	vgain
Xvgain_1		60	60	0	60	vgain
Xvgain_8		60	60	0	60	vgain
Xvgain_32		60	60	0	60	vgain
Xvgain_2		60	60	0	60	vgain
Xvgain_2		60	60	0	60	vgain
Xvgain_2		60	60	0	60	vgain
Xswitch_1		60	60	60	0	switch
Xswitch_1		60	60	60	0	switch
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
XinputI_1		70	60	iin
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvadd_1		60	60	60	60	60	0	60	vadd
Xvtoi_28		0	60	0	vtoi
Xmm_0		0	0	60	60	0	0	0	60	mm
Xmm_0		0	0	60	60	0	0	0	60	mm
XinputV_0		72	60	vin
XinputV_0		72	60	vin
XinputV_2		70	60	vin
XinputV_32		71	60	vin
XinputV_35		68	60	vin
XinputV_23		65	60	vin
XinputV_27		67	60	vin
XinputV_32		71	60	vin
XinputV_1		72	60	vin
XinputV_12		62	60	vin
XinputV_13		69	60	vin
XinputV_1		72	60	vin
XinputV_1		72	60	vin
XinputV_77		71	60	vin
XinputV_1		72	60	vin
XinputV_1		72	60	vin
XinputV_8		66	40	vin
XinputV_1		72	60	vin
XinputV_1		72	60	vin
XinputV_1		72	60	vin
XinputV_1		72	60	vin
Xitov_22		0	0	0	itov
Xitov_8		0	60	60	itov
Xitov_27		60	0	0	itov
Xitov_3		60	0	60	itov
Xitov_9		60	0	60	itov
Xitov_29		60	0	60	itov
Xitov_2		60	0	60	itov
Xitov_17		60	60	0	itov
Xitov_14		0	60	60	itov
Xitov_14		0	60	60	itov
Xitov_29		60	0	60	itov
Xitov_14		0	60	60	itov
Xitov_23		60	0	0	itov
Xitov_0		0	60	60	itov
Xitov_17		60	60	0	itov
Xitov_3		60	0	60	itov
Xitov_11		0	40	0	itov
