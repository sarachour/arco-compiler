
*@input UTF
Iin_UTF_24		79	0	DC	1.
*
*constant value 0.
Vcst23		78	0	DC	0.
*
*constant value 2.5
Vcst22		77	0	DC	2.5
*
*constant value 2.0015
Vcst21		76	0	DC	2.0015
*
*@input umodif
Iin_umodif_20		76	0	DC	1.
*
*@input V
Iin_V_19		75	0	DC	1.
*
*@output U
*@args 74,V
*
*@input VTF
Vin_VTF_17		73	0	DC	1.
*
*constant value 156.25
Icst16		72	0	DC	156.25
*
*@input IPTG
Iin_IPTG_15		71	0	DC	1.
*
*@input V_0
Vin_V_0_14		70	0	DC	1.
*
*constant value 0.01
Vcst13		69	0	DC	0.01
*
*@output umodif
*@args 68,I
*
*@input U_0
Vin_U_0_11		67	0	DC	1.
*
*@output UTF
*@args 67,I
*
*constant value 250.
Vcst9		66	0	DC	250.
*
*@input U
Iin_U_8		65	0	DC	1.
*
*constant value 15.6
Icst7		64	0	DC	15.6
*
*@output V
*@args 63,V
*
*constant value 1.
Vcst5		62	0	DC	1.
*
*@input V
Vin_V_4		61	0	DC	1.
*
*constant value -0.1
Vcst3		60	0	DC	-0.1
*
*constant value 2.9618e-05
Icst2		59	0	DC	2.9618e-05
*
*@output VTF
*@args 58,I
*
*@input Km
Iin_Km_0		57	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_5		48	39	33	7	vgain
Xswitch_0		27	46	21	17	switch
XinputI_1		79	27	iin
XinputI_1		79	27	iin
XinputI_2		59	21	iin
XinputI_7		76	53	iin
XinputI_14		75	11	iin
XinputI_32		72	15	iin
XinputI_24		57	52	iin
XinputI_42		64	42	iin
XinputI_7		76	53	iin
XoutputV_0		44	74	vout
XoutputV_8		5	63	vout
Xvadd_1		32	32	3	40	0	44	35	vadd
Xvadd_32		32	7	32	1	0	5	54	vadd
Xihill_1		15	11	19	52	0	56	ihill
Xihill_6		42	53	39	52	0	56	ihill
XinputV_45		60	9	vin
XinputV_43		69	40	vin
XinputV_40		67	35	vin
XinputV_13		76	46	vin
XinputV_12		66	48	vin
XinputV_46		73	33	vin
XinputV_33		62	39	vin
XinputV_0		70	54	vin
XinputV_37		61	1	vin
XinputV_1		78	32	vin
XinputV_48		77	19	vin
Xitov_14		27	9	3	itov
XoutputI_1		17	68	iout
XoutputI_7		56	67	iout
XoutputI_7		56	67	iout
