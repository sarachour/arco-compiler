EXAMPLE PSpice
*
* ## Dependencies
*
.INCLUDE math/basic.subckt
*
* ## Structure
*
VIN1 1 0 DC 3
VIN2 2 0 DC 5
* plus side of vin1 and vin2
XVMul 1 2 3 VOUT vaddmul

*
* ## Analysis and Plotting
*
.OP
*.TF V(3,0) VIN
*.DC VIN 0 20 2
*.PRINT DC V(1,2) V(2,4) I(VMEAS)
*.PLOT DC V(1,2) V(2,4)
*.PLOT DC I(VMEAS)
.END
