* AD734 SPICE Macro-model
* Description: Amplifier 
* Generic Desc: Bipolar, Multiplier, 4 Quad
* Developed by: AAG / PMI
* Revision History: 08/10/2012 - Updated to new header style
* 2.0 (04/1992) - Removed input signal current compensation: GX1,GY1,GZ1
*		- Added Isy vs. Vsy
* Copyright 1992, 2012 by Analog Devices.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
*
* END Notes

* Node assignments
*             X1
*             |  X2
*             |  |  UO
*             |  |  |  U1
*             |  |  |  |  U2
*             |  |  |  |  |  Y1
*             |  |  |  |  |  |  Y2
*             |  |  |  |  |  |  |  VN
*             |  |  |  |  |  |  |  |   ER
*             |  |  |  |  |  |  |  |   |  Z2
*             |  |  |  |  |  |  |  |   |  |  Z1
*             |  |  |  |  |  |  |  |   |  |  |  W
*             |  |  |  |  |  |  |  |   |  |  |  |  DD
*             |  |  |  |  |  |  |  |   |  |  |  |  |  VP
*             |  |  |  |  |  |  |  |   |  |  |  |  |  |
.SUBCKT AD734 10 11 49 50 51 20 21 200 58 31 30 77 54 100
*
EREF 300 0 POLY(2) 100 0 200 0 (0,0.5,0.5)
*
* X INPUT STAGE & POLE AT 40 MHz
*
CINX 10 11 2E-12
IBX1 10 0 DC 50E-9
IBX2 11 0 DC 50E-9
EOSX 12 10 POLY(1) 18 300 15E-3 1
RX1 12 13 25E3
RX2 13 11 25E3
*
GX1 300 14 12 11 1E-6
RX3 14 300 9.995E5
CX1 14 300 3.9809E-15
VX1 100 15 DC 3.1875
DX1 14 15 DX
VX2 16 200 DC 3.1875
DX2 16 14 DX
*
* X INPUT STAGE COMMON-MODE REJECTION AND ZERO 40 kHz
*
ECMX 17 300 13 300 56.234
RCMX1 17 18 1E6
CCMX 17 18 3.9789E-12
RCMX2 18 300 1
*
* Y INPUT STAGE & POLE AT 40 MHz
*
CINY 20 21 2E-12
IBY1 20 0 DC 50E-9
IBY2 21 0 DC 50E-9
EOSY 22 20 POLY(1) 28 300 10E-3 1
RY1 22 23 25E3
RY2 23 21 25E3
*
GY1 300 24 22 21 1E-6
RY3 24 300 9.995E5
CY1 24 300 3.9809E-15
VY1 100 25 DC 3.1875
DY1 24 25 DX
VY2 26 200 DC 3.1875
DY2 26 24 DX
*
* Y INPUT STAGE COMMON-MODE REJECTION AND ZERO 80 kHz
*
ECMY 27 300 23 300 56.234
RCMY1 27 28 1E6
CCMY 27 28 1.9895E-12
RCMY2 28 300 1
*
* Z INPUT STAGE & POLE AT 40 MHz
*
CINZ 30 31 2E-12
IBZ1 30 0 DC 50E-9
IBZ2 31 0 DC 50E-9
EOSZ 32 30 POLY(1) 38 300 20E-3 1
RZ1 32 33 25E3
RZ2 33 31 25E3
*
GZ1 300 34 32 31 1E-6
RZ3 34 300 1E6
CZ1 34 300 3.9789E-15
VZ1 100 35 DC 3.1875
DZ1 34 35 DX
VZ2 36 200 DC 3.1875
DZ2 36 34 DX
*
* Z INPUT STAGE COMMON-MODE REJECTION AND ZERO 40 kHz
*
ECMZ 37 300 33 300 56.234
RCMZ1 37 38 1E6
CCMZ 37 38 3.9789E-12
RCMZ2 38 300 1
*
* DENOMINATOR CONTROL & INTERNAL REFERENCE
*
QU1 100 49 50 QNU
RU1 50 51 28E3
*
VU 100 52
QU2 52 0 53 QNU
RU2 53 54 0.001
IU 53 200 DC 10E-6
FU1 300 55 VU 1.01
RU3 55 300 1E6
*
VR1 57 200 DC 8
QR 59 57 58 QPU
RR 57 58 1E5
VR2 59 200
FU4 300 56 VR2 1
RU4 56 300 28E3
*
EU 60 300 POLY(3) 50 51 55 300 56 300 (0,1.0101,1,1.0101)
RU5 60 300 1E6
*
* 250 MHz MULTIPLIER CORE
*
EXY 46 300 POLY(2) 14 300 24 300 (0,0,0,0,1)
RXY 46 300 1E6
GXY 300 47 46 300 1
GU 47 300 POLY(2) 60 300 47 300 (0,0,0,0,1)
RU 47 300 1E12
CU 47 300 6.65E-9
EW 48 300 POLY(2) 47 300 34 300 (0,1,-1)
RW 48 300 1E6
*
* OUTPUT AMP BUFFER
*
GW 64 300 48 300 1
QW1 100 0 61 QNW
QW2 200 0 62 QPW
QW3 63 62 64 QNW
QW4 65 61 64 QPW
RW1 100 63 1
RW2 65 200 1
IW1 100 62 DC 100E-6
IW2 61 200 DC 100E-6
VW1 100 66 DC 10
DW1 66 63 DX
VW2 67 200 DC 10
DW2 65 67 DX
*
* OUTPUT AMP GAIN STAGE
*
GW1 300 68 100 63 1
GW2 68 300 65 200 1
RW3 68 300 1.38E3
CW1 68 300 19E-9
VW3 100 69 DC 3.8
DW3 68 69 DX
VW4 70 200 DC 3.8
DW4 70 68 DX
*
* TRANSIENT SUPPLY CURRENT COMPENSATION
*
DCC1 80 100 DX
GCC 0 80 48 300 1
DCC2 0 80 DX
DEE1 81 0 DX
GEE 81 0 300 48 1
DEE2 200 81 DX
*
* POLE AT 17.5 MHz
*
GW3 300 71 68 300 1E-6
RW4 71 300 1E6
CW2 71 300 9.0946E-15
*
IDC 100 200 DC 4.0125E-3
RDC1 100 78 3.2E3
RDC2 78 200 3.2E3
DO1 100 72 DX
GO1 72 200 76 71 25E-3
DO2 200 72 DY
DO3 100 73 DX
GO2 73 200 71 76 25E-3
DO4 200 73 DY
VSC1 74 76 DC 0.4
DSC1 71 74 DX
VSC2 76 75 DC 0.4
DSC2 75 71 DX
GO3 76 100 100 71 25E-3
GO4 200 76 71 200 25E-3
RO1 100 76 40
RO2 76 200 40
LO 76 77 100E-9
*
* MODELS USED
*
.MODEL QNU NPN (BF=100 IS=1E-16)
.MODEL QPU PNP (BF=100 IS=1E-16)
.MODEL QNW NPN (BF=1E9 IS=1E-15)
.MODEL QPW PNP (BF=1E9 IS=1E-15)
.MODEL DX D(IS=1E-15)
.MODEL DY D(IS=1E-15 BV=50)
.ENDS AD734


