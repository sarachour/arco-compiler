
*@input A
Vin_A_2		9	0	DC	1.
*
*@output C
*@args 8,V
*
*constant value 1.
Vcst0		7	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
XoutputV_0		5	8	vout
Xvadd2_2		1	3	5	vadd2
XinputV_8		7	1	vin
XinputV_4		9	3	vin
