
*@input TRLacL
Vin_TRLacL_39		103	0	DC	1.
*
*constant value 0.3010299956
Vcst38		102	0	DC	0.3010299956
*
*constant value 1.
Vcst37		102	0	DC	1.
*
*@input TRTetR
Vin_TRTetR_36		102	0	DC	1.
*
*@input clp
Iin_clp_35		101	0	DC	1.
*
*@input clm
Vin_clm_34		101	0	DC	1.
*
*constant value -0.004
Vcst33		100	0	DC	-0.004
*
*@input TetRp
Iin_TetRp_32		100	0	DC	1.
*
*constant value 0.
Icst31		99	0	DC	0.
*
*@input clp_0
Vin_clp_0_30		99	0	DC	1.
*
*constant value 0.
Vcst29		99	0	DC	0.
*
*@input LacLm_0
Vin_LacLm_0_28		98	0	DC	1.
*
*@output clp
*@args 98,V
*
*@output clm
*@args 98,V
*
*@output TetRm
*@args 98,V
*
*@output LacLm
*@args 98,V
*
*@output LacLp
*@args 98,V
*
*@output TetRp
*@args 97,V
*
*@input TRclp
Iin_TRclp_21		96	0	DC	1.
*
*constant value 0.0005
Icst20		95	0	DC	0.0005
*
*@input TetRp_0
Vin_TetRp_0_19		94	0	DC	1.
*
*@input KM
Iin_KM_18		94	0	DC	1.
*
*@input TRLacL
Iin_TRLacL_17		93	0	DC	1.
*
*constant value -0.1
Vcst16		93	0	DC	-0.1
*
*@input LacLm
Vin_LacLm_15		92	0	DC	1.
*
*@output TRLacL
*@args 92,I
*
*@output TRTetR
*@args 92,I
*
*@output TRclp
*@args 91,I
*
*constant value 752.57498916
Vcst11		91	0	DC	752.57498916
*
*constant value 0.4995
Icst10		90	0	DC	0.4995
*
*constant value 2.
Vcst9		90	0	DC	2.
*
*@input TetRm
Vin_TetRm_8		89	0	DC	1.
*
*@input TetRm_0
Vin_TetRm_0_7		88	0	DC	1.
*
*@input LacLp_0
Vin_LacLp_0_6		87	0	DC	1.
*
*constant value 0.00132877123795
Vcst5		86	0	DC	0.00132877123795
*
*constant value -250.
Vcst4		86	0	DC	-250.
*
*@input clm_0
Vin_clm_0_3		85	0	DC	1.
*
*@input TRclp
Vin_TRclp_2		85	0	DC	1.
*
*constant value 1.5051499783
Vcst1		84	0	DC	1.5051499783
*
*@input LacLp
Iin_LacLp_0		83	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_10		82	82	82	82	vgain
Xvgain_1		82	82	82	82	vgain
Xvgain_4		82	82	82	82	vgain
Xvgain_4		82	82	82	82	vgain
Xvgain_0		82	82	82	82	vgain
Xvgain_1		82	82	82	82	vgain
XinputI_7		83	82	iin
XinputI_48		96	82	iin
XinputI_4		100	82	iin
XinputI_32		95	57	iin
XinputI_15		101	82	iin
XinputI_8		90	12	iin
XinputI_2		94	82	iin
XoutputV_4		82	98	vout
Xvadd_32		82	82	82	82	0	82	82	vadd
Xvadd_33		82	82	82	82	0	82	79	vadd
Xvadd_29		82	82	82	82	0	82	30	vadd
Xihill_4		12	82	82	82	0	82	ihill
Xihill_2		12	82	82	82	0	82	ihill
Xihill_5		12	82	82	82	0	82	ihill
XinputV_5		91	82	vin
XinputV_38		86	82	vin
XinputV_4		88	79	vin
XinputV_48		102	82	vin
XinputV_48		102	82	vin
XinputV_16		101	82	vin
XinputV_48		102	82	vin
XinputV_22		103	82	vin
XinputV_9		87	79	vin
XinputV_1		86	82	vin
XinputV_8		93	82	vin
XinputV_30		94	30	vin
XinputV_2		90	82	vin
XinputV_5		91	82	vin
Xitov_1		82	82	82	itov
Xiadd_18		57	82	82	82	82	iadd
Xiadd_10		57	82	82	82	82	iadd
XoutputI_0		82	92	iout
