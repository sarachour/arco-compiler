
*constant value 0.00132877123795
Vcst38		132	0	DC	0.00132877123795
*
*@output clp
*@args 131,V
*
*@output TetRm
*@args 131,V
*
*constant value 1.
Vcst35		130	0	DC	1.
*
*constant value -0.0005
Icst34		129	0	DC	-0.0005
*
*constant value 1.5051499783
Vcst33		129	0	DC	1.5051499783
*
*constant value 0.0005
Icst32		128	0	DC	0.0005
*
*@input TetRm_0
Vin_TetRm_0_31		128	0	DC	1.
*
*@input TetRp
Iin_TetRp_30		128	0	DC	1.
*
*constant value -0.1
Vcst29		128	0	DC	-0.1
*
*@output TetRp
*@args 127,V
*
*@input KM
Iin_KM_27		126	0	DC	1.
*
*@output TRTetR
*@args 126,I
*
*@input TRLacL
Vin_TRLacL_25		126	0	DC	1.
*
*@output LacLm
*@args 126,V
*
*constant value 0.
Vcst23		126	0	DC	0.
*
*@input LacLm_0
Vin_LacLm_0_22		126	0	DC	1.
*
*@output TRLacL
*@args 125,I
*
*@input clp
Iin_clp_20		124	0	DC	1.
*
*@input clp_0
Vin_clp_0_19		124	0	DC	1.
*
*constant value 2.
Vcst18		123	0	DC	2.
*
*constant value 0.
Icst17		122	0	DC	0.
*
*@input TetRp_0
Vin_TetRp_0_16		121	0	DC	1.
*
*constant value 0.4995
Icst15		120	0	DC	0.4995
*
*constant value 0.004
Vcst14		119	0	DC	0.004
*
*@output LacLp
*@args 118,V
*
*@output TRclp
*@args 117,I
*
*@input clm
Vin_clm_11		116	0	DC	1.
*
*@input TRclp
Vin_TRclp_10		115	0	DC	1.
*
*constant value 752.57498916
Vcst9		115	0	DC	752.57498916
*
*@input TetRm
Vin_TetRm_8		114	0	DC	1.
*
*@input LacLm
Vin_LacLm_7		114	0	DC	1.
*
*@input LacLp_0
Vin_LacLp_0_6		114	0	DC	1.
*
*@input TRTetR
Iin_TRTetR_5		113	0	DC	1.
*
*constant value -250.
Vcst4		112	0	DC	-250.
*
*@output clm
*@args 111,V
*
*@input clm_0
Vin_clm_0_2		110	0	DC	1.
*
*@input LacLp
Iin_LacLp_1		109	0	DC	1.
*
*constant value 0.3010299956
Vcst0		108	0	DC	0.3010299956
*
*
*
* === Connectivity Schem ==== 
Xvgain_5		19	104	1	104	vgain
Xvgain_25		104	104	19	74	vgain
Xvgain_6		104	19	104	24	vgain
Xvgain_35		19	104	80	59	vgain
Xvgain_2		104	19	104	106	vgain
XinputI_11		113	3	iin
XinputI_35		124	30	iin
XinputI_33		128	36	iin
XinputI_20		122	13	iin
XinputI_46		120	87	iin
XinputI_48		128	82	iin
XinputI_44		126	29	iin
XinputI_15		129	49	iin
XinputI_48		128	82	iin
XoutputV_8		78	131	vout
XoutputV_7		78	111	vout
XoutputV_0		99	126	vout
XoutputV_0		99	126	vout
XoutputV_8		78	131	vout
XoutputV_4		32	131	vout
Xvadd_28		104	104	104	104	0	78	104	vadd
Xvadd_28		104	104	104	104	0	78	104	vadd
Xvadd_24		74	104	104	40	0	99	104	vadd
Xvadd_33		104	104	24	104	0	99	104	vadd
Xvadd_1		59	104	104	40	0	78	46	vadd
Xvadd_2		106	104	104	40	0	32	104	vadd
Xihill_2		87	30	58	29	0	70	ihill
Xihill_5		87	82	58	29	0	51	ihill
Xihill_0		87	82	58	29	0	66	ihill
XinputV_48		132	104	vin
XinputV_1		129	104	vin
XinputV_2		119	104	vin
XinputV_39		115	1	vin
XinputV_48		132	104	vin
XinputV_25		116	104	vin
XinputV_48		132	104	vin
XinputV_48		132	104	vin
XinputV_19		108	40	vin
XinputV_48		132	104	vin
XinputV_42		123	58	vin
XinputV_1		129	104	vin
XinputV_48		132	104	vin
XinputV_1		129	104	vin
XinputV_31		130	19	vin
XinputV_1		129	104	vin
XinputV_1		129	104	vin
XinputV_40		121	46	vin
XinputV_36		114	80	vin
XinputV_48		132	104	vin
XinputV_1		129	104	vin
Xitov_2		3	104	104	itov
Xiadd_15		70	36	13	13	53	iadd
Xiadd_28		36	51	13	13	77	iadd
Xiadd_0		13	66	13	49	77	iadd
XoutputI_3		53	117	iout
XoutputI_8		77	126	iout
XoutputI_8		77	126	iout
