
*constant value 0.3010299956
Vcst41		65	0	DC	0.3010299956
*
*constant value 30.1029995664
Icst40		65	0	DC	30.1029995664
*
*constant value 0.0005
Icst32		65	0	DC	0.0005
*
*@input TetRm_0
Vin_TetRm_0_30		65	0	DC	1.
*
*constant value 10
Vcst28		65	0	DC	10.
*
*@input LacLp_0
Vin_LacLp_0_25		65	0	DC	1.
*
*constant value 0
Icst19		64	0	DC	0.
*
*@input clp_0
Vin_clp_0_16		63	0	DC	1.
*
*constant value 0.4995
Icst13		61	0	DC	0.4995
*
*constant value 30.1029995664
Vcst11		59	0	DC	30.1029995664
*
*constant value 10
Icst10		58	0	DC	10.
*
*constant value 0
Vcst9		57	0	DC	0.
*
*@input TetRp_0
Vin_TetRp_0_8		56	0	DC	1.
*
*@input LacLm_0
Vin_LacLm_0_7		56	0	DC	1.
*
*constant value 2
Vcst4		54	0	DC	2.
*
*@input clm_0
Vin_clm_0_3		53	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
XinputI_25		65	21	iin
XinputI_0		65	51	iin
XinputI_14		65	51	iin
XinputI_4		65	51	iin
XinputI_0		65	51	iin
Xvadd_0		51	51	51	51	0	0	51	vadd
Xvadd_0		51	51	51	51	0	0	51	vadd
Xvadd_0		51	51	51	51	0	0	51	vadd
Xvadd_0		51	51	51	51	0	0	51	vadd
Xvadd_6		51	13	51	0	0	0	51	vadd
Xvadd_3		51	51	51	0	0	0	3	vadd
Xihill_1		51	0	51	0	0	19	ihill
Xihill_0		51	0	51	0	0	35	ihill
Xihill_4		51	0	51	0	0	35	ihill
XinputV_0		65	51	vin
XinputV_0		65	51	vin
XinputV_28		65	51	vin
XinputV_123		65	51	vin
XinputV_104		65	51	vin
XinputV_1		65	51	vin
XinputV_0		65	51	vin
XinputV_117		65	51	vin
XinputV_28		65	51	vin
XinputV_116		65	3	vin
XinputV_58		65	51	vin
Xitov_2		0	51	51	itov
Xitov_9		0	51	51	itov
Xitov_17		21	0	51	itov
Xitov_26		51	0	51	itov
Xitov_10		0	51	13	itov
Xitov_9		0	51	51	itov
Xiadd_21		51	19	51	51	0	iadd
Xiadd_0		51	35	51	51	0	iadd
Xiadd_0		51	35	51	51	0	iadd
