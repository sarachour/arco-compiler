
*@input IPTG
Iin_IPTG_28		39	0	DC	1.
*
*@input U_0
Vin_U_0_27		39	0	DC	1.
*
*constant value 0
Vcst26		39	0	DC	0.
*
*constant value 15.6
Icst22		38	0	DC	15.6
*
*constant value 2.9618e-05
Icst19		36	0	DC	2.9618e-05
*
*constant value 10
Vcst18		36	0	DC	10.
*
*constant value 10
Icst17		36	0	DC	10.
*
*constant value 156.25
Icst13		36	0	DC	156.25
*
*constant value 2.0015
Vcst9		35	0	DC	2.0015
*
*constant value 0.01
Vcst7		33	0	DC	0.01
*
*@input V_0
Vin_V_0_5		31	0	DC	1.
*
*constant value 1
Vcst3		29	0	DC	1.
*
*constant value 2.5
Vcst2		29	0	DC	2.5
*
*
*
* === Connectivity Schem ==== 
Xswitch_5		26	13	21	0	switch
XinputI_29		39	23	iin
XinputI_0		39	18	iin
XinputI_17		39	21	iin
XinputI_12		39	26	iin
XinputI_0		39	18	iin
Xvadd_0		26	26	26	11	0	0	26	vadd
Xvadd_0		26	26	26	11	0	0	26	vadd
Xihill_6		23	0	5	0	0	0	ihill
Xihill_5		18	0	13	0	0	0	ihill
XinputV_89		36	5	vin
XinputV_119		36	26	vin
XinputV_72		36	11	vin
XinputV_83		39	26	vin
XinputV_25		36	26	vin
XinputV_113		39	26	vin
XinputV_0		35	13	vin
XinputV_0		35	13	vin
Xitov_26		0	26	26	itov
Xitov_22		18	0	26	itov
