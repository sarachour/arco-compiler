
*@input ES_0
Iin_ES_0_6		22	0	DC	1.
*
*@output S
*@args 21,I
*
*@output E
*@args 20,I
*
*constant value 1.
Icst3		19	0	DC	1.
*
*@output ES
*@args 18,I
*
*constant value 0.15
Icst1		17	0	DC	0.15
*
*constant value 0.11
Icst0		16	0	DC	0.11
*
*
*
* === Connectivity Schem ==== 
XinputI_2		17	10	iin
XinputI_46		19	3	iin
XinputI_4		22	12	iin
XinputI_47		16	8	iin
Xmm_0		8	10	3	3	14	4	6	12	mm
XoutputI_7		14	18	iout
XoutputI_0		4	21	iout
XoutputI_9		6	20	iout
