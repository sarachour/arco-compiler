
*@output C
*@args 9,I
*
*@input A
Iin_A_0		8	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
XinputI_0		8	7	iin
Ximul2_3		1	7	3	imul2
XoutputI_2		3	9	iout
XcopyI_1		7	1	icopy
