
*@input R_0
Vin_R_0_92		108	0	DC	1.
*
*@input MA_0
Vin_MA_0_90		108	0	DC	1.
*
*@input DR_0
Vin_DR_0_85		108	0	DC	1.
*
*constant value -10
Vcst84		108	0	DC	-10.
*
*constant value 0.01
Icst80		108	0	DC	0.01
*
*@input DRp_0
Vin_DRp_0_75		108	0	DC	1.
*
*constant value 0.0008
Vcst74		108	0	DC	0.0008
*
*constant value 0
Vcst71		108	0	DC	0.
*
*constant value 10
Vcst68		108	0	DC	10.
*
*@input C_0
Vin_C_0_65		108	0	DC	1.
*
*constant value 0.2
Icst60		108	0	DC	0.2
*
*constant value -100
Vcst59		108	0	DC	-100.
*
*constant value 250
Vcst56		108	0	DC	250.
*
*constant value -100
Icst54		107	0	DC	-100.
*
*constant value 0
Icst49		106	0	DC	0.
*
*constant value 2500
Vcst48		106	0	DC	2500.
*
*constant value -1
Vcst47		106	0	DC	-1.
*
*constant value 0.2
Vcst46		106	0	DC	0.2
*
*@input MR_0
Vin_MR_0_45		106	0	DC	1.
*
*constant value 0.010101010101
Icst43		106	0	DC	0.010101010101
*
*constant value 0.00200400801603
Icst39		105	0	DC	0.00200400801603
*
*constant value 12.5
Vcst37		105	0	DC	12.5
*
*constant value 10
Icst36		105	0	DC	10.
*
*constant value 50
Vcst35		104	0	DC	50.
*
*constant value 50
Icst34		104	0	DC	50.
*
*constant value 0.04
Vcst30		104	0	DC	0.04
*
*constant value 1
Icst25		102	0	DC	1.
*
*@input DAp_0
Vin_DAp_0_19		99	0	DC	1.
*
*constant value 0.0204081632653
Icst18		99	0	DC	0.0204081632653
*
*@input A_0
Vin_A_0_15		98	0	DC	1.
*
*constant value 1
Vcst11		96	0	DC	1.
*
*@input DA_0
Vin_DA_0_10		95	0	DC	1.
*
*constant value 0.004
Vcst7		94	0	DC	0.004
*
*constant value 49
Icst4		92	0	DC	49.
*
*
*
* === Connectivity Schem ==== 
Xvgain_2		59	89	0	89	vgain
Xvgain_37		59	89	0	89	vgain
Xvgain_3		89	89	0	89	vgain
Xvgain_31		89	89	0	89	vgain
Xvgain_38		89	89	0	71	vgain
Xvgain_4		89	89	0	89	vgain
Xvgain_7		89	89	0	48	vgain
Xvgain_36		89	89	0	0	vgain
Xswitch_0		7	89	89	0	switch
Xswitch_2		89	89	89	0	switch
Xswitch_9		89	89	89	0	switch
Xswitch_5		89	89	89	0	switch
XinputI_21		108	7	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
XinputI_1		105	89	iin
XinputI_22		108	80	iin
XinputI_0		108	89	iin
XinputI_0		108	89	iin
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvadd_6		89	71	89	89	0	0	89	vadd
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvadd_15		89	48	89	89	0	0	85	vadd
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvadd_0		89	89	89	89	89	0	89	vadd
Xvtoi_28		0	89	0	vtoi
Xmm_0		0	0	89	89	0	0	0	89	mm
Xmm_0		0	0	89	89	0	0	0	89	mm
XinputV_79		108	41	vin
XinputV_56		108	89	vin
XinputV_19		108	83	vin
XinputV_54		106	59	vin
XinputV_38		108	65	vin
XinputV_68		104	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_20		108	89	vin
XinputV_0		108	89	vin
XinputV_5		106	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_24		106	89	vin
XinputV_12		108	85	vin
XinputV_23		108	89	vin
XinputV_41		108	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_0		108	89	vin
XinputV_13		108	89	vin
Xitov_13		0	41	0	itov
Xitov_28		89	0	89	itov
Xitov_28		89	0	89	itov
Xitov_16		0	83	89	itov
Xitov_23		0	65	89	itov
Xitov_21		0	89	89	itov
Xitov_18		0	89	89	itov
Xitov_15		89	0	0	itov
Xitov_12		0	0	0	itov
Xitov_18		0	89	89	itov
Xitov_8		80	0	0	itov
Xitov_14		0	0	0	itov
Xitov_28		89	0	89	itov
Xitov_2		89	0	0	itov
Xitov_9		0	89	89	itov
