
*constant value 1
Vcst30		72	0	DC	1.
*
*@input TetRp_0
Vin_TetRp_0_29		72	0	DC	1.
*
*constant value 0.4995
Icst28		72	0	DC	0.4995
*
*constant value 2
Vcst27		72	0	DC	2.
*
*constant value 30.1029995664
Icst26		71	0	DC	30.1029995664
*
*@input LacLm_0
Vin_LacLm_0_25		70	0	DC	1.
*
*constant value 0
Icst23		69	0	DC	0.
*
*constant value 30.1029995664
Vcst21		68	0	DC	30.1029995664
*
*@input LacLp_0
Vin_LacLp_0_20		68	0	DC	1.
*
*constant value 0.0005
Icst18		67	0	DC	0.0005
*
*constant value 0.004
Vcst17		66	0	DC	0.004
*
*constant value 250
Vcst13		66	0	DC	250.
*
*constant value 0.3010299956
Vcst11		66	0	DC	0.3010299956
*
*constant value 752.57498916
Vcst9		66	0	DC	752.57498916
*
*constant value 0
Vcst8		65	0	DC	0.
*
*@input clp_0
Vin_clp_0_7		64	0	DC	1.
*
*constant value 1.5051499783
Vcst6		64	0	DC	1.5051499783
*
*@input clm_0
Vin_clm_0_4		63	0	DC	1.
*
*@input TetRm_0
Vin_TetRm_0_2		62	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_1		61	61	0	61	vgain
Xvgain_2		61	40	0	61	vgain
Xvgain_0		61	61	0	58	vgain
Xvgain_15		61	61	0	61	vgain
XinputI_1		72	61	iin
XinputI_0		69	61	iin
XinputI_31		67	45	iin
XinputI_1		72	61	iin
Xvadd_1		61	61	61	61	0	0	61	vadd
Xvadd_1		61	61	61	61	0	0	61	vadd
Xvadd_7		61	58	61	61	0	0	61	vadd
Xvadd_3		61	13	61	0	0	0	17	vadd
Xvadd_1		61	61	61	61	0	0	61	vadd
Xvadd_1		61	61	61	61	0	0	61	vadd
Xihill_7		61	0	61	0	0	29	ihill
Xihill_1		61	0	61	0	0	19	ihill
Xihill_6		61	0	61	0	0	22	ihill
XinputV_0		66	61	vin
XinputV_2		66	40	vin
XinputV_6		64	61	vin
XinputV_3		72	61	vin
XinputV_0		66	61	vin
XinputV_6		64	61	vin
XinputV_3		72	61	vin
XinputV_1		72	61	vin
XinputV_46		64	17	vin
XinputV_1		72	61	vin
XinputV_1		72	61	vin
XinputV_1		72	61	vin
XinputV_1		72	61	vin
XinputV_1		72	61	vin
XinputV_14		68	61	vin
Xitov_9		61	0	13	itov
Xitov_17		0	61	61	itov
Xiadd_0		45	29	61	61	0	iadd
Xiadd_16		45	19	61	61	0	iadd
Xiadd_24		45	22	61	61	0	iadd
