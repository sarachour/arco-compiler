
*@input DAp_0
Vin_DAp_0_81		88	0	DC	1.
*
*constant value 50
Vcst80		88	0	DC	50.
*
*@input C_0
Vin_C_0_75		88	0	DC	1.
*
*constant value 10
Vcst73		88	0	DC	10.
*
*constant value 0.5
Icst71		88	0	DC	0.5
*
*constant value 0.0008
Vcst64		88	0	DC	0.0008
*
*constant value 0
Vcst62		88	0	DC	0.
*
*constant value 10
Icst60		88	0	DC	10.
*
*@input MR_0
Vin_MR_0_58		87	0	DC	1.
*
*constant value 0
Icst53		87	0	DC	0.
*
*constant value 0.2
Vcst51		86	0	DC	0.2
*
*@input DR_0
Vin_DR_0_49		86	0	DC	1.
*
*constant value 1
Icst44		84	0	DC	1.
*
*@input MA_0
Vin_MA_0_43		84	0	DC	1.
*
*constant value 500
Vcst35		83	0	DC	500.
*
*@input DRp_0
Vin_DRp_0_34		82	0	DC	1.
*
*constant value 0.01
Vcst31		82	0	DC	0.01
*
*constant value 50
Icst30		82	0	DC	50.
*
*@input A_0
Vin_A_0_25		82	0	DC	1.
*
*constant value -10
Vcst20		80	0	DC	-10.
*
*@input R_0
Vin_R_0_17		78	0	DC	1.
*
*constant value 1
Vcst14		77	0	DC	1.
*
*constant value -100
Vcst10		76	0	DC	-100.
*
*@input DA_0
Vin_DA_0_9		75	0	DC	1.
*
*constant value 100
Icst0		72	0	DC	100.
*
*
*
* === Connectivity Schem ==== 
Xvgain_10		0	71	0	0	vgain
XinputI_28		88	71	iin
XinputI_0		88	71	iin
XinputI_0		88	71	iin
XinputI_0		88	71	iin
XinputI_0		88	71	iin
XinputI_0		88	71	iin
Xvadd_11		71	71	71	0	0	0	71	vadd
Xvadd_10		30	71	71	0	0	0	13	vadd
Xvadd_0		71	71	71	71	63	0	71	vadd
Xvadd_0		71	71	71	71	63	0	71	vadd
Xvadd_31		47	63	54	0	0	0	28	vadd
Xvadd_0		71	71	71	71	63	0	71	vadd
Xvadd_0		71	71	71	71	63	0	71	vadd
Xvadd_0		71	71	71	71	63	0	71	vadd
Xvtoi_0		0	71	0	vtoi
Xvtoi_0		0	71	0	vtoi
Xvtoi_28		0	71	0	vtoi
Xmm_0		0	0	71	71	0	0	0	71	mm
Xmm_0		0	0	71	71	0	0	0	71	mm
XinputV_40		87	71	vin
XinputV_0		88	71	vin
XinputV_57		88	71	vin
XinputV_61		82	71	vin
XinputV_14		88	71	vin
XinputV_0		88	71	vin
XinputV_0		88	71	vin
XinputV_6		88	71	vin
XinputV_0		88	71	vin
XinputV_20		88	71	vin
XinputV_106		88	13	vin
XinputV_85		88	71	vin
XinputV_0		88	71	vin
XinputV_42		83	71	vin
XinputV_60		82	28	vin
XinputV_67		86	71	vin
XinputV_0		88	71	vin
XinputV_7		86	71	vin
XinputV_91		83	71	vin
Xitov_8		71	71	71	itov
Xitov_2		71	71	71	itov
Xitov_27		0	71	0	itov
Xitov_1		71	71	71	itov
Xitov_26		0	71	71	itov
Xitov_10		71	0	0	itov
Xitov_24		0	71	71	itov
Xitov_13		71	71	30	itov
Xitov_1		71	71	71	itov
Xitov_1		71	71	71	itov
Xitov_18		0	0	0	itov
Xitov_19		0	71	0	itov
Xitov_26		0	71	71	itov
Xitov_12		0	71	47	itov
Xitov_4		0	71	54	itov
Xitov_8		71	71	71	itov
Xitov_0		71	71	71	itov
Xitov_0		71	71	71	itov
Xitov_3		71	0	71	itov
Xitov_1		71	71	71	itov
Xitov_2		71	71	71	itov
Xitov_13		71	71	30	itov
Xitov_27		0	71	0	itov
Xitov_6		71	71	71	itov
Xitov_6		71	71	71	itov
Xitov_0		71	71	71	itov
