
*@output UTF
*@args 60,I
*
*@input V
Vin_V_12		59	0	DC	1.
*
*constant value 15.6
Icst11		58	0	DC	15.6
*
*@input IPTG
Vin_IPTG_10		57	0	DC	1.
*
*@input U
Vin_U_9		56	0	DC	1.
*
*constant value 156.25
Icst8		55	0	DC	156.25
*
*@input umodif
Iin_umodif_7		54	0	DC	1.
*
*@output umodif
*@args 53,V
*
*constant value 1.
Icst5		52	0	DC	1.
*
*constant value 1.
Vcst4		51	0	DC	1.
*
*@output VTF
*@args 50,I
*
*constant value -2.0015
Vcst2		50	0	DC	-2.0015
*
*constant value 2.5
Vcst1		49	0	DC	2.5
*
*constant value 33763.2520764
Icst0		48	0	DC	33763.2520764
*
*
*
* === Connectivity Schem ==== 
Xvgain_19		43	11	43	1	vgain
Xvgain_38		43	29	23	27	vgain
Xvgain_20		43	9	43	3	vgain
Xswitch_2		31	20	25	5	switch
XinputI_2		48	31	iin
XinputI_47		52	15	iin
XinputI_29		58	7	iin
XinputI_34		54	21	iin
XinputI_30		55	33	iin
XoutputV_2		27	53	vout
Xihill_0		33	15	20	46	0	44	ihill
Xvtoi_4		43	1	25	vtoi
Xvtoi_3		3	43	46	vtoi
Xigenebind_2		21	15	7	16	igenebind
XinputV_25		57	11	vin
XinputV_8		56	23	vin
XinputV_1		50	20	vin
XinputV_13		51	43	vin
XinputV_14		59	9	vin
Xitov_4		5	43	29	itov
XoutputI_0		16	50	iout
XoutputI_7		44	60	iout
