EXAMPLE PSpice
*
* ## Dependencies
*
.INCLUDE libs/basic.subckt
*
* ## Structure
*
VIN1 c1 0 DC 1
VIN2 c2 0 DC 2
VSIN1 sin1 0 DC SIN(0V 5V 100Hz) 



rin sin1 in 0
*rout sin1 out 0
xcmp sin1 out 0 vvderiv
*xcmp sin1 out 0 vvinteg
*xcmp in1 in2 0 out vadd

*
* ## Analysis and Plotting
*
.control
	set stime=1us
	set etime=0.01s

	op
	tran $stime $etime 
	
	gnuplot out-trans:in tran.V(in)
	gnuplot out-trans:out tran.V(out)
.endc


.END




*.TF V(out,0) VSIN1
*.PRINT DC V(out,0)
*.SENS V(out,0)
*.DISPLAY
