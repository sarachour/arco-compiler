
*@input B
Vin_B_4		19	0	DC	#
*
*@input A
Vin_A_3		18	0	DC	#
*
*@input A
Vin_A_2		17	0	DC	#
*
*@output C
*@args 16 V
*
*@input A
Vin_A_0		15	0	DC	#
*
*
*
* === Connectivity Schem ====
XoutputV_1		11	16	vout
Xvadd2_3		7	13	11	vadd2
XinputV_2		15	1	vin
XinputV_3		18	9	vin
XinputV_8		17	5	vin
XinputV_1		19	3	vin
Xvmul2_1		1	9	13	vmul2
Xvmul2_3		3	5	7	vmul2
