
*@output U
*@args 58,I
*
*@output V
*@args 57,I
*
*constant value 156.25
Icst19		56	0	DC	156.25
*
*@input VTF
Iin_VTF_18		55	0	DC	1.
*
*@input U_0
Iin_U_0_17		55	0	DC	1.
*
*@input V_0
Iin_V_0_16		54	0	DC	1.
*
*@input UTF
Iin_UTF_15		54	0	DC	1.
*
*constant value 0.001
Icst14		53	0	DC	0.001
*
*@input U
Iin_U_13		52	0	DC	1.
*
*constant value 0.
Icst12		51	0	DC	0.
*
*@output UTF
*@args 51,I
*
*@output VTF
*@args 50,I
*
*@input umodif
Iin_umodif_9		49	0	DC	1.
*
*constant value 15.6
Icst8		48	0	DC	15.6
*
*@input IPTG
Iin_IPTG_7		47	0	DC	1.
*
*constant value 2.0015
Icst6		46	0	DC	2.0015
*
*@output umodif
*@args 45,I
*
*constant value -1.
Icst4		44	0	DC	-1.
*
*@input V
Iin_V_3		43	0	DC	1.
*
*constant value 1.
Icst2		42	0	DC	1.
*
*constant value -2.5
Icst1		42	0	DC	-2.5
*
*constant value 2.9618e-05
Icst0		41	0	DC	2.9618e-05
*
*
*
* === Connectivity Schem ==== 
Xswitch_9		40	23	23	26	switch
Xadd4_19		33	33	24	3	0	add4
Xmult4_1		12	23	26	23	38	mult4
XinputI_10		43	24	iin
XinputI_36		44	3	iin
XinputI_8		51	33	iin
XinputI_4		56	7	iin
XinputI_14		55	18	iin
XinputI_0		54	18	iin
XinputI_15		55	36	iin
XinputI_1		48	7	iin
XinputI_34		42	23	iin
XinputI_24		49	26	iin
XinputI_25		52	12	iin
XinputI_12		46	23	iin
XinputI_5		42	23	iin
XinputI_2		47	40	iin
Xstateful_14		18	18	27	0	stateful
Xinh_bind_4		26	7	23	23	29	inhbind
XoutputI_5		27	58	iout
XoutputI_4		29	51	iout
XoutputI_3		38	45	iout
