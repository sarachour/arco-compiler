
*@input E_0
Vin_E_0_28		33	0	DC	1.
*
*constant value 25.25
Icst26		33	0	DC	25.25
*
*constant value 0.0190476190476
Vcst24		33	0	DC	0.0190476190476
*
*@output P
Vout_P_19		33	0	DC	1.
*
*@input ES_0
Vin_ES_0_17		32	0	DC	1.
*
*constant value 1
Vcst15		32	0	DC	1.
*
*constant value 0.00172786177106
Vcst14		32	0	DC	0.00172786177106
*
*constant value 0.00126823081801
Vcst10		31	0	DC	0.00126823081801
*
*constant value 0
Vcst9		31	0	DC	0.
*
*@input S_0
Vin_S_0_7		30	0	DC	1.
*
*@input P_0
Vin_P_0_6		30	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_28		15	25	0	25	vgain
Xvgain_20		25	0	0	25	vgain
Xvgain_14		0	25	0	25	vgain
Xvgain_18		15	25	0	25	vgain
XinputI_0		33	23	iin
XoutputV_0		33	0	vout
Xvadd_0		25	25	25	0	0	20	25	vadd
Xvadd_0		25	25	25	0	0	20	25	vadd
Xvadd_0		25	25	25	0	0	20	25	vadd
Xvadd_0		25	25	25	0	0	20	25	vadd
XinputV_61		33	25	vin
XinputV_5		32	15	vin
XinputV_122		33	25	vin
XinputV_0		33	25	vin
XinputV_7		31	25	vin
XinputV_122		33	25	vin
XinputV_0		33	25	vin
XinputV_34		32	25	vin
XinputV_0		33	25	vin
Xitov_3		23	0	25	itov
