
*@input S
Vin_S_18		32	0	DC	1.
*
*constant value 0.760456273764
Vcst17		32	0	DC	0.760456273764
*
*@input E
Vin_E_16		31	0	DC	1.
*
*constant value -0.317057704502
Vcst15		30	0	DC	-0.317057704502
*
*constant value 0.
Vcst14		30	0	DC	0.
*
*@input P_0
Vin_P_0_13		29	0	DC	1.
*
*@output ES
*@args 29,V
*
*@output P
*@args 29,V
*
*@input ES
Iin_ES_10		28	0	DC	1.
*
*constant value 1.
Vcst9		27	0	DC	1.
*
*@output E
*@args 27,V
*
*@output S
*@args 26,V
*
*constant value 0.655737704918
Vcst6		26	0	DC	0.655737704918
*
*@input ES
Vin_ES_5		26	0	DC	1.
*
*constant value -4.7619047619
Vcst4		25	0	DC	-4.7619047619
*
*@input E_0
Vin_E_0_3		25	0	DC	1.
*
*@input S_0
Vin_S_0_2		25	0	DC	1.
*
*@input ES_0
Vin_ES_0_1		24	0	DC	1.
*
*constant value 2.525
Vcst0		23	0	DC	2.525
*
*
*
* === Connectivity Schem ==== 
Xvgain_0		23	23	23	23	vgain
Xvgain_0		23	23	23	23	vgain
XinputI_25		28	23	iin
XoutputV_0		23	29	vout
XoutputV_0		23	29	vout
Xvadd_1		23	23	23	23	0	23	23	vaddgain
XinputV_17		27	23	vin
XinputV_4		25	23	vin
XinputV_27		23	23	vin
XinputV_13		32	23	vin
XinputV_0		32	23	vin
XinputV_9		30	23	vin
XinputV_1		30	23	vin
XinputV_0		32	23	vin
Xitov_0		23	23	23	itov
Xitov_0		23	23	23	itov
