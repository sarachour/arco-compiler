
*@output UTF
*@args 64,I
*
*@output VTF
*@args 63,I
*
*constant value 156.25
Icst11		63	0	DC	156.25
*
*@input umodif
Iin_umodif_10		62	0	DC	1.
*
*@input V
Iin_V_9		61	0	DC	1.
*
*constant value 1.
Vcst8		61	0	DC	1.
*
*@output umodif
*@args 60,V
*
*constant value 33763.2520764
Icst6		59	0	DC	33763.2520764
*
*constant value 2.5
Vcst5		58	0	DC	2.5
*
*constant value -2.0015
Vcst4		57	0	DC	-2.0015
*
*@input U
Vin_U_3		56	0	DC	1.
*
*@input IPTG
Vin_IPTG_2		55	0	DC	1.
*
*@input Km
Iin_Km_1		55	0	DC	1.
*
*constant value 15.6
Icst0		54	0	DC	15.6
*
*
*
* === Connectivity Schem ==== 
Xvgain_12		42	48	42	23	vgain
Xvgain_10		42	48	42	12	vgain
Xvgain_34		42	48	42	43	vgain
Xswitch_0		27	42	21	23	switch
Xswitch_2		27	42	42	23	switch
XinputI_41		59	27	iin
XinputI_14		61	51	iin
XinputI_23		55	51	iin
XinputI_15		63	51	iin
XoutputV_0		43	60	vout
Xihill_6		51	51	42	51	0	52	ihill
Xvtoi_9		23	42	21	vtoi
Xvtoi_2		12	42	42	vtoi
Xvtoi_1		43	42	42	vtoi
Xvtoi_13		12	42	42	vtoi
XinputV_43		55	48	vin
XinputV_25		61	42	vin
XinputV_19		56	42	vin
XinputV_25		61	42	vin
XinputV_0		58	42	vin
Xitov_3		23	42	48	itov
Xitov_3		23	42	48	itov
Xitov_2		23	42	48	itov
XoutputI_0		52	64	iout
