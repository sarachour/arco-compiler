
*@output P
*@args 63,V
*
*@output E
*@args 63,V
*
*constant value 578.75
Vcst14		63	0	DC	578.75
*
*@input S
Vin_S_13		62	0	DC	1.
*
*@input E
Vin_E_12		61	0	DC	1.
*
*@output ES
*@args 60,V
*
*constant value 0.0190476190476
Vcst10		60	0	DC	0.0190476190476
*
*constant value 0.00126823081801
Vcst9		59	0	DC	0.00126823081801
*
*constant value 1.
Vcst8		58	0	DC	1.
*
*@input P_0
Vin_P_0_7		57	0	DC	1.
*
*@input ES_0
Vin_ES_0_6		56	0	DC	1.
*
*constant value 631.25
Vcst5		55	0	DC	631.25
*
*@output S
*@args 54,V
*
*@input E_0
Vin_E_0_3		53	0	DC	1.
*
*@input ES
Vin_ES_2		52	0	DC	1.
*
*@input S_0
Vin_S_0_1		51	0	DC	1.
*
*constant value 0.
Vcst0		50	0	DC	0.
*
*
*
* === Connectivity Schem ==== 
Xvgain_4		45	47	16	1	vgain
Xvgain_14		38	12	44	49	vgain
Xvgain_21		38	12	44	49	vgain
Xvgain_35		12	38	44	27	vgain
XoutputV_10		3	60	vout
XoutputV_60		38	63	vout
XoutputV_60		38	63	vout
XoutputV_1		35	63	vout
Xvadd_33		31	1	24	44	0	3	25	vadd
Xvadd_4		24	49	24	16	0	38	38	vadd
Xvadd_4		24	49	24	16	0	38	38	vadd
Xvadd_9		27	24	24	0	0	35	16	vadd
XinputV_4		59	47	vin
XinputV_110		61	45	vin
XinputV_117		56	25	vin
XinputV_47		55	38	vin
XinputV_120		63	38	vin
XinputV_108		50	24	vin
XinputV_59		62	16	vin
XinputV_0		51	38	vin
XinputV_76		58	12	vin
XinputV_91		52	44	vin
XinputV_120		63	38	vin
XinputV_75		57	16	vin
XinputV_120		63	38	vin
Xitov_3		0	24	31	itov
