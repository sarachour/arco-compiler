* AD834 SPICE Macro-model
* Description: Amplifier 
* Generic Desc: Multiplier, 4 Quad
* Developed by: PN
* Rev 0: Jul 17, 2014
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* Node assignments
*             Y1
*             |  Y2
*             |  | -Vs
*             |  |  |  W2   
*             |  |  |  | W1  
*             |  |  |  |  | +Vs  
*             |  |  |  |  |  |  X1  
*             |  |  |  |  |  |  | X2
*             |  |  |  |  |  |  |  |   
.SUBCKT AD834 Y1 Y2 50 W2 W1 99 X1 X2

*X differential input stage

R19 X2 5 1e-006 
R18 X1 4 1e-006

*Bias current
I2 5 98  4.5e-005 
I1 4 98  4.5e-005

*Input Clamp
D14 4 11 Diode
V26 11 5  1.3 
D13 20 4 Diode
V23 5 20  1.3 

*CMR
R2 6 5 12500 
R1 4 6 12500 
E17 4 3 10 98 1
C2 9 10 3.1e-011
R4 9 10 3830 
R3 98 10 1 
E2 9 98 6 98 1

*input offset X
V1 3 7  0.0005 

*Input X Amplifier
R29 5 12 1000 
R28 7 21 1000 
R27 21 Xout 1000 
R13 12 98 1000 
G7 Xout 98 13 98 1
C3 13 98 2.65258e-010
R5 13 98 100000 
G3 13 98 21 12 1

V13 45 50  1 
D5 45 44 Diode
V11 99 43 1 
D4 Xout 43 Diode

*Distortion 
G12 Xout1 98 Xout 98 3e-005
L1 23 98 1.5915e-005
R21 Xout1 23 1100 
xA6 Xout1 98 A6_OPEN_3 A6_OPEN_4 A6_OPEN_5 A6_OPEN_6 22 98 POLYSourceA6
.SUBCKT POLYSourceA6 1 2 3 4 5 6 7 8
E1 7 8 POLY(3) (1,2) (3,4) (5,6) 0 0 0 0 1 0 0 0 0 0  0 0 0 0 0
R0 1 2 1e15
R1 3 4 1e15
R2 5 6 1e15
R3 5 0 1e15
R4 3 0 1e15
R5 1 0 1e15
.ENDS

xA3 22 98 Xout 98 A3_OPEN_5 A3_OPEN_6 Xout2 98 POLYSourceA3
.SUBCKT POLYSourceA3 1 2 3 4 5 6 7 8
E1 7 8 POLY(3) (1,2) (3,4) (5,6) 0 1 1 0 0 0 0 0 0 0  0 0 0 0 0
R0 1 2 1e15
R1 3 4 1e15
R2 5 6 1e15
R3 5 0 1e15
R4 3 0 1e15
R5 1 0 1e15
.ENDS

V6 99 41 1 
D2 Xout2 41 Diode
V10 42 50 1 
D3 42 Xout2 Diode

*Y Differential input stage

R26 Y2 15 1e-006 
R25 Y1 14 1e-006 

*Bias current
I5 15 98  4.5e-005
I4 14 98 4.5e-005 

*Input clamp
D7 14 1 Diode
V20 1 15 1.3 
D6 18 14 Diode
V16 15 18  1.3 

*CMR
E12 14 37 28 98 1
C1 27 28 3.1e-011
R10 27 28 3830 
R9 98 28 1 
E9 27 98 26 98 1
R8 26 15 12500 
R7 14 26 12500 

*Input Offset Y
V8 37 16  0.0005

*Input Y Amplifier
R33 15 30 1000 
R32 16 29 1000 
R31 29 Yout 1000 
R30 30 98 1000 
G8 Yout 98 31 98 1
C4 31 98 2.65258e-010
R11 31 98 100000 
G6 31 98 29 30 1

V24 99 49 1 
D11 Yout 49 Diode
V18 46 50 1 
D8 46 Yout Diode

*Distortion
G13 Yout1 98 Yout 98 2e-005
L2 25 98 1.5915e-005
R20 Yout1 25 1100 

xA8 Yout1 98 A8_OPEN_3 A8_OPEN_4 A8_OPEN_5 A8_OPEN_6 24 98 POLYSourceA8
.SUBCKT POLYSourceA8 1 2 3 4 5 6 7 8
E1 7 8 POLY(3) (1,2) (3,4) (5,6) 0 0 0 0 1 0 0 0 0 0  0 0 0 0 0
R0 1 2 1e15
R1 3 4 1e15
R2 5 6 1e15
R3 5 0 1e15
R4 3 0 1e15
R5 1 0 1e15
.ENDS

xA7 24 98 Yout 98 A7_OPEN_5 A7_OPEN_6 Yout2 98 POLYSourceA7
.SUBCKT POLYSourceA7 1 2 3 4 5 6 7 8
E1 7 8 POLY(3) (1,2) (3,4) (5,6) 0 1 1 0 0 0 0 0 0 0  0 0 0 0 0
R0 1 2 1e15
R1 3 4 1e15
R2 5 6 1e15
R3 5 0 1e15
R4 3 0 1e15
R5 1 0 1e15
.ENDS

V21 99 48  1 
D10 Yout2 48 Diode
V19 47 50 1 
D9 47 Yout2 Diode

*Multiplier Core
xA1 Xout2 98 Yout2 98 A1_OPEN_5 A1_OPEN_6 xy_out 98 POLYSourceA1
.SUBCKT POLYSourceA1 1 2 3 4 5 6 7 8
E1 7 8 POLY(3) (1,2) (3,4) (5,6) 0 0 0 0 0 1 0 0 0 0  0 0 0 0 0
R0 1 2 1e15
R1 3 4 1e15
R2 5 6 1e15
R3 5 0 1e15
R4 3 0 1e15
R5 1 0 1e15
.ENDS

*Noise
V4 40 98  0.6 
R6 38 98 15 
D1 40 39 DNoise
E3 17 xy_out 38 39 0.0037

*Output Amplifier
E15 out 98 35 34 1
R22 98 33 1000 
R35 out 32 1000 
R16 17 32 1000 
R12 33 98 1000 
C6 35 34 2e-010
R34 35 34 100000
G14 35 34 32 33 1
G9 W1 W2 out 98 0.004

*Differential Offset Output Current
I17 W1 W2  2e-005 

*Standing Output Current
I11 W1 98 0.0085 
I10 W2 98  0.0085
 
*Quiescent Current
I16 99 98  0.011 
I15 50 98  0.028 

*diode model
.model Diode  D
.model DNoise  D
+ (
+  KF=3.4e-019
+ )
 
.ENDS AD834

