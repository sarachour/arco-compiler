
*@output S
*@args 27,I
*
*@output ES
*@args 27,I
*
*@output P
*@args 27,I
*
*@output E
*@args 26,I
*
*constant value 1.01
Icst9		26	0	DC	1.01
*
*@input P_0
Iin_P_0_8		25	0	DC	1.
*
*@input E
Iin_E_7		25	0	DC	1.
*
*constant value 1.
Icst6		24	0	DC	1.
*
*@input ES
Iin_ES_5		23	0	DC	1.
*
*@input S_0
Iin_S_0_4		23	0	DC	1.
*
*@input ES_0
Iin_ES_0_3		23	0	DC	1.
*
*@input E_0
Iin_E_0_2		22	0	DC	1.
*
*@input S
Iin_S_1		22	0	DC	1.
*
*constant value 0.01
Icst0		21	0	DC	0.01
*
*
*
* === Connectivity Schem ==== 
Xmult4_1		20	20	20	20	20	mult4
Xmult4_17		20	20	20	20	20	mult4
XinputI_49		26	20	iin
XinputI_5		23	20	iin
XinputI_25		22	20	iin
XinputI_48		25	20	iin
XinputI_1		23	20	iin
Xstateful_4		20	20	9	0	stateful
XoutputI_1		9	27	iout
