
*@output MA
*@args 136,V
*
*constant value 50.
Vcst43		136	0	DC	50.
*
*@output MR
*@args 136,V
*
*@output DR
*@args 135,V
*
*@input C
Vin_C_40		134	0	DC	1.
*
*@output C
*@args 133,V
*
*@input DA
Vin_DA_38		132	0	DC	1.
*
*@input MA
Vin_MA_37		132	0	DC	1.
*
*@output DA
*@args 132,V
*
*@input DR_0
Vin_DR_0_35		132	0	DC	1.
*
*@input C_0
Vin_C_0_34		131	0	DC	1.
*
*@input DAp_0
Vin_DAp_0_33		130	0	DC	1.
*
*@input A
Vin_A_32		129	0	DC	1.
*
*constant value -8e-06
Vcst31		128	0	DC	-8e-06
*
*@input MA_0
Vin_MA_0_30		128	0	DC	1.
*
*@input DA_0
Vin_DA_0_29		128	0	DC	1.
*
*@output DRp
*@args 128,V
*
*constant value -0.004
Vcst27		127	0	DC	-0.004
*
*constant value 0.
Vcst26		127	0	DC	0.
*
*@input A_0
Vin_A_0_25		126	0	DC	1.
*
*@output DAp
*@args 126,V
*
*constant value -10000.
Vcst23		125	0	DC	-10000.
*
*@input R_0
Vin_R_0_22		124	0	DC	1.
*
*@input MR_0
Vin_MR_0_21		124	0	DC	1.
*
*@input MR
Iin_MR_20		123	0	DC	1.
*
*@input MR
Vin_MR_19		123	0	DC	1.
*
*@input DR
Vin_DR_18		122	0	DC	1.
*
*constant value 1.
Vcst17		121	0	DC	1.
*
*constant value 250.
Vcst16		120	0	DC	250.
*
*constant value 8e-05
Vcst15		120	0	DC	8e-05
*
*@output A
*@args 119,V
*
*@output R
*@args 118,V
*
*@input DA
Iin_DA_12		117	0	DC	1.
*
*constant value -100.
Icst11		116	0	DC	-100.
*
*constant value 125000.
Vcst10		116	0	DC	125000.
*
*@input R
Vin_R_9		116	0	DC	1.
*
*constant value 0.004
Vcst8		116	0	DC	0.004
*
*constant value 0.02
Vcst7		115	0	DC	0.02
*
*@input DRp
Vin_DRp_6		114	0	DC	1.
*
*@input DRp_0
Vin_DRp_0_5		113	0	DC	1.
*
*constant value 0.1
Icst4		112	0	DC	0.1
*
*constant value 500.
Vcst3		111	0	DC	500.
*
*constant value 1000.
Vcst2		110	0	DC	1000.
*
*@input DAp
Vin_DAp_1		109	0	DC	1.
*
*@input DRp
Iin_DRp_0		108	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_2		107	107	107	107	vgain
Xvgain_20		107	10	107	8	vgain
Xvgain_3		107	47	107	53	vgain
Xvgain_0		107	107	107	107	vgain
Xvgain_38		107	107	107	107	vgain
Xvgain_11		107	107	107	107	vgain
Xvgain_38		107	107	107	107	vgain
Xvgain_0		107	107	107	107	vgain
Xvgain_38		107	107	107	107	vgain
Xvgain_34		107	107	107	89	vgain
Xvgain_0		107	107	107	107	vgain
XinputI_9		123	107	iin
XinputI_3		117	107	iin
XinputI_22		116	81	iin
XinputI_6		108	107	iin
XinputI_23		112	50	iin
XoutputV_58		107	133	vout
XoutputV_72		107	136	vout
XoutputV_13		74	118	vout
XoutputV_26		107	136	vout
XoutputV_72		107	136	vout
XoutputV_34		107	135	vout
XoutputV_72		107	136	vout
XoutputV_72		107	136	vout
XoutputV_72		107	136	vout
Xvadd_32		107	107	107	107	0	107	107	vadd
Xvadd_5		107	107	8	107	0	107	107	vadd
Xvadd_14		107	107	53	107	0	74	14	vadd
Xvadd_32		107	107	107	107	0	107	107	vadd
Xvadd_25		107	12	107	107	29	0	0	vadd
Xvadd_33		107	29	107	107	0	107	56	vadd
Xvadd_32		107	107	107	107	0	107	107	vadd
Xvadd_10		107	89	107	107	0	107	76	vadd
Xvadd_32		107	107	107	107	0	107	107	vadd
Xvadd_32		107	107	107	107	0	107	107	vadd
XinputV_103		131	107	vin
XinputV_54		127	10	vin
XinputV_123		136	107	vin
XinputV_122		132	107	vin
XinputV_123		136	107	vin
XinputV_121		115	47	vin
XinputV_113		120	107	vin
XinputV_120		134	107	vin
XinputV_71		124	14	vin
XinputV_98		111	107	vin
XinputV_123		136	107	vin
XinputV_123		136	107	vin
XinputV_115		109	107	vin
XinputV_117		132	107	vin
XinputV_84		128	107	vin
XinputV_38		121	107	vin
XinputV_60		125	107	vin
XinputV_20		132	107	vin
XinputV_4		129	107	vin
XinputV_117		132	107	vin
XinputV_122		132	107	vin
XinputV_3		126	56	vin
XinputV_122		132	107	vin
XinputV_122		132	107	vin
XinputV_122		132	107	vin
XinputV_5		110	58	vin
XinputV_47		130	76	vin
XinputV_122		132	107	vin
XinputV_122		132	107	vin
XinputV_122		132	107	vin
XinputV_122		132	107	vin
Xitov_24		107	107	107	itov
Xitov_24		107	107	107	itov
Xitov_16		81	107	12	itov
Xitov_24		107	107	107	itov
Xitov_17		107	58	107	itov
Xitov_28		50	107	107	itov
Xitov_7		107	107	107	itov
