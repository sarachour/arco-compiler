
*@output E
*@args 57,V
*
*constant value 25.25
Vcst17		57	0	DC	25.25
*
*@input S
Vin_S_16		56	0	DC	1.
*
*@input E
Vin_E_15		55	0	DC	1.
*
*@output P
*@args 54,V
*
*@input E_0
Vin_E_0_13		54	0	DC	1.
*
*constant value 2.1
Icst12		53	0	DC	2.1
*
*@input P_0
Vin_P_0_11		53	0	DC	1.
*
*@input ES
Iin_ES_10		52	0	DC	1.
*
*constant value 0.00126823081801
Vcst9		52	0	DC	0.00126823081801
*
*constant value 23.15
Vcst8		52	0	DC	23.15
*
*constant value 1.
Vcst7		51	0	DC	1.
*
*constant value 631.25
Vcst6		51	0	DC	631.25
*
*@output S
*@args 50,V
*
*@input ES
Vin_ES_4		49	0	DC	1.
*
*@output ES
*@args 48,V
*
*@input S_0
Vin_S_0_2		48	0	DC	1.
*
*@input ES_0
Vin_ES_0_1		47	0	DC	1.
*
*constant value 0.
Vcst0		46	0	DC	0.
*
*
*
* === Connectivity Schem ==== 
Xvgain_37		0	0	37	31	vgain
Xvgain_7		1	45	37	3	vgain
Xvgain_38		37	23	45	37	vgain
XinputI_47		52	33	iin
XinputI_48		53	28	iin
XoutputV_53		5	48	vout
XoutputV_72		45	57	vout
XoutputV_0		7	50	vout
XoutputV_72		45	57	vout
Xvadd_23		31	3	37	45	0	5	45	vadd
Xvadd_32		37	37	37	37	0	45	45	vadd
Xvadd_14		37	9	37	37	0	7	45	vadd
Xvadd_32		37	37	37	37	0	45	45	vadd
XinputV_26		55	1	vin
XinputV_122		57	45	vin
XinputV_122		57	45	vin
XinputV_122		57	45	vin
XinputV_123		51	37	vin
XinputV_99		49	45	vin
XinputV_9		51	23	vin
XinputV_122		57	45	vin
XinputV_123		51	37	vin
XinputV_80		56	37	vin
XinputV_122		57	45	vin
XinputV_122		57	45	vin
XinputV_122		57	45	vin
Xitov_27		33	45	9	itov
Xitov_28		28	45	37	itov
