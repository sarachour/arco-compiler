
*@output E
*@args 22,V
*
*@output S
*@args 21,V
*
*constant value 0.11
Vcst5		20	0	DC	0.11
*
*constant value 0.15
Vcst4		19	0	DC	0.15
*
*@input ES_0
Vin_ES_0_3		18	0	DC	1.
*
*constant value 1.
Icst2		18	0	DC	1.
*
*@output ES
*@args 17,V
*
*@input ES
Iin_ES_0		16	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
XinputI_48		18	13	iin
XinputI_48		18	13	iin
XoutputV_73		14	17	vout
XoutputV_71		3	21	vout
XoutputV_64		1	22	vout
Xmm_0		9	7	13	13	14	1	3	5	mm
XinputV_52		18	5	vin
XinputV_7		20	7	vin
XinputV_75		19	9	vin
