
*constant value 0.
Icst9		29	0	DC	0.
*
*@input ES_0
Vin_ES_0_8		28	0	DC	1.
*
*@output E
*@args 28,V
*
*@output ES
*@args 27,V
*
*constant value 0.2
Icst5		26	0	DC	0.2
*
*@input Q
Iin_Q_4		25	0	DC	1.
*
*@output S
*@args 24,V
*
*constant value 0.11
Vcst2		24	0	DC	0.11
*
*constant value 0.15
Vcst1		23	0	DC	0.15
*
*constant value 20.3
Icst0		22	0	DC	20.3
*
*
*
* === Connectivity Schem ==== 
XinputI_2		25	19	iin
XinputI_0		29	13	iin
XinputI_0		29	13	iin
XinputI_1		26	17	iin
XoutputV_1		21	28	iout
XoutputV_0		3	24	iout
XoutputV_1		21	28	iout
Xmm_0		14	14	7	17	21	3	21	15	mm
XinputV_0		24	14	iin
XinputV_0		24	14	iin
XinputV_3		28	15	iin
Xiadd_1		13	1	7	iadd
Xigain_1		13	19	1	iadd
