
*constant value 23.15
Icst14		30	0	DC	23.15
*
*@output P
Vout_P_13		30	0	DC	1.
*
*constant value 2.1
Icst12		29	0	DC	2.1
*
*constant value 0
Vcst9		28	0	DC	0.
*
*@input P_0
Vin_P_0_8		28	0	DC	1.
*
*constant value 0.00126823081801
Vcst7		28	0	DC	0.00126823081801
*
*@input S_0
Vin_S_0_5		27	0	DC	1.
*
*constant value 25.25
Vcst4		26	0	DC	25.25
*
*@input ES_0
Vin_ES_0_3		25	0	DC	1.
*
*@input E_0
Vin_E_0_1		24	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_2		0	0	23	23	vgain
Xvgain_8		0	23	0	23	vgain
XinputI_1		30	22	iin
XinputI_1		30	22	iin
XoutputV_16		30	0	vout
Xvadd_1		23	23	23	23	0	20	23	vadd
Xvadd_1		23	23	23	23	0	20	23	vadd
Xvadd_1		23	23	23	23	0	20	23	vadd
Xvadd_1		23	23	23	23	0	20	23	vadd
XinputV_97		26	10	vin
XinputV_3		24	23	vin
XinputV_14		27	23	vin
XinputV_8		28	23	vin
XinputV_1		28	23	vin
XinputV_1		28	23	vin
XinputV_1		28	23	vin
Xitov_12		0	10	23	itov
Xitov_23		22	0	23	itov
Xitov_10		22	0	23	itov
