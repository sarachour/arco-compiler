EXAMPLE PSpice
*
* ## Dependencies
*
.INCLUDE math/basic.subckt
*
* ## Structure
*
VIN1 1 0 DC 10
VIN2 2 0 DC 10

x1 1 2 3 vadd
x2 1 3 4 vadd

*
* ## Analysis and Plotting
*
.OP
.END
