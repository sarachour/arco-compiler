
*@output BH3
*@args 514,I
*
*constant value 0.333333333333
Icst177		513	0	DC	0.333333333333
*
*@output BiPT
*@args 513,V
*
*@output WFS1
*@args 513,V
*
*constant value -5.
Icst174		513	0	DC	-5.
*
*@input CHOP
Vin_CHOP_173		513	0	DC	1.
*
*@input Gamma
Iin_Gamma_172		513	0	DC	1.
*
*@output mWFS1
*@args 513,V
*
*@input BH3T
Iin_BH3T_170		513	0	DC	1.
*
*@input mXbp1u_0
Vin_mXbp1u_0_169		513	0	DC	1.
*
*constant value 1.2
Vcst168		513	0	DC	1.2
*
*constant value 0.1
Vcst167		513	0	DC	0.1
*
*@input IRE1
Vin_IRE1_166		513	0	DC	1.
*
*@input WFS1_0
Vin_WFS1_0_165		513	0	DC	1.
*
*@output BH3T
*@args 512,V
*
*@input PERKA
Iin_PERKA_163		512	0	DC	1.
*
*constant value 1.6e-05
Vcst162		512	0	DC	1.6e-05
*
*constant value -0.5
Vcst161		512	0	DC	-0.5
*
*@input ATF4_0
Vin_ATF4_0_160		512	0	DC	1.
*
*@output ATF6
*@args 511,V
*
*constant value -1.05263157895
Icst158		511	0	DC	-1.05263157895
*
*constant value -30.
Vcst157		510	0	DC	-30.
*
*constant value 0.0002
Icst156		510	0	DC	0.0002
*
*@input BAXmBCL2_0
Vin_BAXmBCL2_0_155		510	0	DC	1.
*
*@input BiRE1_0
Vin_BiRE1_0_154		510	0	DC	1.
*
*@input ATF6p50
Vin_ATF6p50_153		510	0	DC	1.
*
*@input ATF6p50
Iin_ATF6p50_152		510	0	DC	1.
*
*@input ATF6T_0
Vin_ATF6T_0_151		510	0	DC	1.
*
*@input IRE1
Iin_IRE1_150		509	0	DC	1.
*
*constant value 2000.
Vcst149		508	0	DC	2000.
*
*constant value 0.004
Vcst148		507	0	DC	0.004
*
*@input BiPER
Iin_BiPER_147		507	0	DC	1.
*
*@input BCL2T
Vin_BCL2T_146		506	0	DC	1.
*
*@input BiPT
Iin_BiPT_145		506	0	DC	1.
*
*@input ATF6GB_0
Vin_ATF6GB_0_144		506	0	DC	1.
*
*constant value 2.
Vcst143		506	0	DC	2.
*
*constant value 25.
Vcst142		505	0	DC	25.
*
*constant value -25000.
Icst141		504	0	DC	-25000.
*
*@input BiRE1
Iin_BiRE1_140		504	0	DC	1.
*
*constant value 1.
Icst139		504	0	DC	1.
*
*@input BiPER_0
Vin_BiPER_0_138		503	0	DC	1.
*
*constant value 10.
Icst137		502	0	DC	10.
*
*@output BiRE1
*@args 501,V
*
*constant value 2.
Icst135		500	0	DC	2.
*
*@input mXbp1s
Vin_mXbp1s_134		499	0	DC	1.
*
*@output mCHOP
*@args 499,V
*
*@input ATF4
Vin_ATF4_132		498	0	DC	1.
*
*constant value 0.0025
Icst131		498	0	DC	0.0025
*
*@input IRE1A
Vin_IRE1A_130		497	0	DC	1.
*
*@output GADD34
*@args 497,V
*
*constant value 0.25
Vcst128		497	0	DC	0.25
*
*@input mWFS1
Vin_mWFS1_127		496	0	DC	1.
*
*@output BAXm
*@args 496,I
*
*@output mGADD34
*@args 495,V
*
*@input mXbp1s_0
Vin_mXbp1s_0_124		494	0	DC	1.
*
*constant value 0.
Vcst123		494	0	DC	0.
*
*constant value 100.
Vcst122		494	0	DC	100.
*
*constant value 4.
Vcst121		494	0	DC	4.
*
*@input BCL2T
Iin_BCL2T_120		493	0	DC	1.
*
*@input eIF2a
Vin_eIF2a_119		493	0	DC	1.
*
*@output ATF4
*@args 493,V
*
*@input mGADD34_0
Vin_mGADD34_0_117		492	0	DC	1.
*
*@input BAXmT_0
Vin_BAXmT_0_116		491	0	DC	1.
*
*@input spliceRate
Vin_spliceRate_115		491	0	DC	1.
*
*@input fGK
Iin_fGK_114		490	0	DC	1.
*
*@output ATF6GB
*@args 490,V
*
*@output mXbp1s
*@args 490,V
*
*constant value 1000000000.
Vcst111		490	0	DC	1000000000.
*
*@input BiRE1
Vin_BiRE1_110		489	0	DC	1.
*
*constant value -5e-05
Icst109		488	0	DC	-5e-05
*
*@input WFS1
Vin_WFS1_108		487	0	DC	1.
*
*constant value -0.1
Vcst107		487	0	DC	-0.1
*
*@input BH3BCL2
Iin_BH3BCL2_106		487	0	DC	1.
*
*@output IRE1
*@args 487,I
*
*@output BCL2T
*@args 487,V
*
*@input mXbp1u
Vin_mXbp1u_103		487	0	DC	1.
*
*@output fGK
*@args 487,V
*
*@input BiPT
Vin_BiPT_101		486	0	DC	1.
*
*@input BAXmT
Iin_BAXmT_100		486	0	DC	1.
*
*@input ATF6T
Vin_ATF6T_99		485	0	DC	1.
*
*@input BiUFP_0
Vin_BiUFP_0_98		484	0	DC	1.
*
*constant value 3000.
Icst97		484	0	DC	3000.
*
*@input BH3BCL2_0
Vin_BH3BCL2_0_96		484	0	DC	1.
*
*constant value 100.
Icst95		484	0	DC	100.
*
*@output ATF6T
*@args 484,V
*
*constant value 0.5
Vcst93		483	0	DC	0.5
*
*@input ATF4
Iin_ATF4_92		483	0	DC	1.
*
*@output eIF2a
*@args 482,I
*
*@input mUFPT
Vin_mUFPT_90		482	0	DC	1.
*
*@input Xbp1s_0
Vin_Xbp1s_0_89		481	0	DC	1.
*
*constant value 4e-05
Vcst88		480	0	DC	4e-05
*
*@output spliceRate
*@args 479,I
*
*constant value 0.03
Icst86		478	0	DC	0.03
*
*@output BH3BCL2
*@args 478,V
*
*@output PERKA
*@args 477,V
*
*@output BiATF
*@args 476,V
*
*@output BiUFP
*@args 476,V
*
*constant value -1.01
Icst81		475	0	DC	-1.01
*
*@input CHOP
Iin_CHOP_80		475	0	DC	1.
*
*@output mBiPT
*@args 475,V
*
*@input BiATF_0
Vin_BiATF_0_78		475	0	DC	1.
*
*@output ATF6p50
*@args 475,V
*
*@input PERKA
Vin_PERKA_76		475	0	DC	1.
*
*@input mCHOP_0
Vin_mCHOP_0_75		474	0	DC	1.
*
*@output Gamma
*@args 473,I
*
*constant value 0.005
Vcst73		473	0	DC	0.005
*
*constant value -1.02564102564
Icst72		472	0	DC	-1.02564102564
*
*@output UFP
*@args 472,V
*
*@output BiPER
*@args 472,V
*
*constant value 0.66666666667
Icst69		471	0	DC	0.66666666667
*
*constant value -1.
Icst68		470	0	DC	-1.
*
*constant value 0.
Icst67		469	0	DC	0.
*
*constant value 20.
Icst66		468	0	DC	20.
*
*constant value -2.
Vcst65		467	0	DC	-2.
*
*@input BAXm
Vin_BAXm_64		466	0	DC	1.
*
*constant value -4.
Vcst63		465	0	DC	-4.
*
*@input UFPT
Vin_UFPT_62		465	0	DC	1.
*
*constant value -10.
Vcst61		465	0	DC	-10.
*
*constant value 20.5
Vcst60		465	0	DC	20.5
*
*@input GADD34
Vin_GADD34_59		464	0	DC	1.
*
*@input mBiPT
Vin_mBiPT_58		463	0	DC	1.
*
*@input ATF6
Vin_ATF6_57		462	0	DC	1.
*
*@input Xbp1s
Vin_Xbp1s_56		462	0	DC	1.
*
*constant value 1.
Vcst55		461	0	DC	1.
*
*@input BiP
Vin_BiP_54		460	0	DC	1.
*
*constant value -100.
Icst53		460	0	DC	-100.
*
*constant value 4.44444444444e-05
Vcst52		459	0	DC	4.44444444444e-05
*
*@output Xbp1s
*@args 459,V
*
*@input BiPT_0
Vin_BiPT_0_50		458	0	DC	1.
*
*@input PERK
Iin_PERK_49		457	0	DC	1.
*
*constant value -1.05
Icst48		457	0	DC	-1.05
*
*@output BAXmBCL2
*@args 457,V
*
*constant value -1.
Vcst46		457	0	DC	-1.
*
*@output CHOP
*@args 456,V
*
*constant value 0.0004
Vcst44		455	0	DC	0.0004
*
*@input BAXmBCL2
Iin_BAXmBCL2_43		455	0	DC	1.
*
*@output PERK
*@args 454,I
*
*@output BiP
*@args 454,V
*
*constant value -1.11111111111
Icst40		453	0	DC	-1.11111111111
*
*@input BH3T_0
Vin_BH3T_0_39		452	0	DC	1.
*
*@output IRE1A
*@args 451,V
*
*@input CHOP_0
Vin_CHOP_0_37		450	0	DC	1.
*
*constant value 250.
Vcst36		449	0	DC	250.
*
*@input IRE1A_0
Vin_IRE1A_0_35		448	0	DC	1.
*
*@output BAXmT
*@args 448,V
*
*constant value 50.
Vcst33		447	0	DC	50.
*
*@output mXbp1u
*@args 446,V
*
*@input mGADD34
Iin_mGADD34_31		445	0	DC	1.
*
*@input PERK
Vin_PERK_30		445	0	DC	1.
*
*@input UFP
Iin_UFP_29		445	0	DC	1.
*
*@input mCHOP
Vin_mCHOP_28		444	0	DC	1.
*
*@input mWFS1_0
Vin_mWFS1_0_27		443	0	DC	1.
*
*@output UFPT
*@args 442,V
*
*@input ATF6p50_0
Vin_ATF6p50_0_25		442	0	DC	1.
*
*constant value 10.
Vcst24		441	0	DC	10.
*
*@input BH3BCL2
Vin_BH3BCL2_23		440	0	DC	1.
*
*constant value 6.
Icst22		440	0	DC	6.
*
*constant value 0.04
Vcst21		440	0	DC	0.04
*
*@input ATF6GB
Vin_ATF6GB_20		439	0	DC	1.
*
*@input BH3T
Vin_BH3T_19		438	0	DC	1.
*
*constant value -250.
Vcst18		437	0	DC	-250.
*
*@input GADD34_0
Vin_GADD34_0_17		436	0	DC	1.
*
*@input UFPT_0
Vin_UFPT_0_16		435	0	DC	1.
*
*constant value -1000.
Vcst15		434	0	DC	-1000.
*
*constant value -0.0566037735848
Icst14		434	0	DC	-0.0566037735848
*
*@input PERKA_0
Vin_PERKA_0_13		433	0	DC	1.
*
*@input mBiPT_0
Vin_mBiPT_0_12		432	0	DC	1.
*
*@input BCL2
Vin_BCL2_11		431	0	DC	1.
*
*constant value 4.
Icst10		430	0	DC	4.
*
*constant value 500.
Vcst9		430	0	DC	500.
*
*@input BH3
Vin_BH3_8		429	0	DC	1.
*
*@input mGADD34
Vin_mGADD34_7		428	0	DC	1.
*
*@output BCL2
*@args 427,I
*
*@input mBiPT
Iin_mBiPT_5		427	0	DC	1.
*
*constant value -2500.
Vcst4		426	0	DC	-2500.
*
*@input BCL2T_0
Vin_BCL2T_0_3		425	0	DC	1.
*
*@input mCHOP
Iin_mCHOP_2		424	0	DC	1.
*
*@input GADD34
Iin_GADD34_1		423	0	DC	1.
*
*@input mXbp1u
Iin_mXbp1u_0		422	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_13		422	422	422	422	vgain
Xvgain_6		422	422	422	422	vgain
Xvgain_2		422	422	422	422	vgain
Xvgain_6		422	422	422	422	vgain
Xvgain_2		422	422	422	422	vgain
Xvgain_18		422	422	422	422	vgain
Xvgain_34		422	422	422	422	vgain
Xvgain_36		422	422	422	422	vgain
Xvgain_2		422	422	422	422	vgain
Xvgain_36		422	422	422	422	vgain
Xvgain_2		422	422	422	422	vgain
Xvgain_4		422	422	422	422	vgain
Xvgain_30		0	0	422	303	vgain
Xvgain_5		422	340	422	342	vgain
Xvgain_38		422	340	422	422	vgain
Xvgain_13		422	422	422	422	vgain
Xvgain_18		422	422	422	422	vgain
Xvgain_35		422	422	422	422	vgain
Xvgain_37		422	422	422	422	vgain
Xvgain_28		422	422	246	422	vgain
Xvgain_9		327	422	422	422	vgain
Xvgain_7		254	62	327	422	vgain
Xvgain_28		422	422	246	422	vgain
Xvgain_25		422	422	422	9	vgain
Xvgain_16		422	422	422	223	vgain
Xvgain_1		422	422	422	422	vgain
Xvgain_22		422	368	422	422	vgain
Xvgain_3		422	422	422	368	vgain
Xswitch_11		422	422	422	422	switch
Xswitch_4		422	422	422	422	switch
Xswitch_12		422	422	422	422	switch
Xswitch_13		422	422	422	422	switch
Xswitch_12		422	422	422	422	switch
Xswitch_3		422	422	422	422	switch
Xswitch_10		422	422	422	422	switch
Xswitch_1		422	422	422	422	switch
Xswitch_5		422	422	422	422	switch
Xswitch_4		422	422	422	422	switch
Xswitch_4		422	422	422	422	switch
Xswitch_13		422	422	422	422	switch
Xswitch_0		422	422	422	387	switch
Xswitch_1		422	422	422	422	switch
Xswitch_5		422	422	422	422	switch
XinputI_20		500	422	iin
XinputI_34		430	422	iin
XinputI_47		513	422	iin
XinputI_47		513	422	iin
XinputI_47		513	422	iin
XinputI_47		513	422	iin
XinputI_2		483	422	iin
XinputI_10		488	11	iin
XinputI_2		483	422	iin
XinputI_1		511	422	iin
XinputI_1		511	422	iin
XinputI_48		513	422	iin
XinputI_19		513	422	iin
XinputI_24		468	422	iin
XinputI_22		457	422	iin
XinputI_47		513	422	iin
XinputI_4		470	422	iin
XinputI_12		493	97	iin
XinputI_48		513	422	iin
XinputI_42		502	422	iin
XinputI_44		510	422	iin
XinputI_45		504	422	iin
XinputI_43		469	422	iin
XinputI_45		504	422	iin
XinputI_46		510	422	iin
XinputI_44		510	422	iin
XinputI_47		513	422	iin
XinputI_48		513	422	iin
XinputI_45		504	422	iin
XinputI_47		513	422	iin
XinputI_48		513	422	iin
XinputI_46		510	422	iin
XinputI_33		490	422	iin
XinputI_38		424	422	iin
XinputI_47		513	422	iin
XinputI_45		504	422	iin
XinputI_39		509	422	iin
XinputI_48		513	422	iin
XinputI_46		510	422	iin
XinputI_47		513	422	iin
XinputI_36		504	422	iin
XinputI_47		513	422	iin
XinputI_28		472	422	iin
XinputI_48		513	422	iin
XinputI_48		513	422	iin
XinputI_44		510	422	iin
XinputI_48		513	422	iin
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_69		422	476	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_39		422	495	vout
XoutputV_9		422	478	vout
XoutputV_6		41	512	vout
XoutputV_72		422	513	vout
XoutputV_23		422	501	vout
XoutputV_72		422	513	vout
XoutputV_16		422	497	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_69		422	476	vout
XoutputV_0		422	513	vout
XoutputV_15		422	511	vout
XoutputV_0		422	513	vout
XoutputV_9		422	478	vout
XoutputV_14		422	487	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_16		422	497	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_72		422	513	vout
XoutputV_14		422	487	vout
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_33		422	422	422	422	0	422	422	vadd
Xvadd_4		114	422	422	422	0	422	87	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_28		303	422	422	422	0	41	422	vadd
Xvadd_16		422	342	422	422	0	422	19	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_33		422	422	422	422	0	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_15		422	422	422	422	0	422	422	vadd
Xvadd_32		422	422	422	422	422	422	422	vadd
Xvadd_8		422	422	422	422	0	422	422	vadd
Xvadd_0		422	422	422	395	0	422	422	vadd
Xvadd_21		9	422	422	422	246	0	0	vadd
Xvadd_2		422	422	223	422	0	422	422	vadd
Xihill_3		422	422	422	422	0	0	ihill
Xihill_5		422	422	422	422	0	422	ihill
Xihill_5		422	422	422	422	0	422	ihill
Xihill_5		422	422	422	422	0	422	ihill
Xvtoi_27		422	422	422	vtoi
Xvtoi_16		422	166	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xvtoi_13		422	422	422	vtoi
Xvtoi_2		422	346	104	vtoi
Xvtoi_1		422	422	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xvtoi_11		422	422	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xvtoi_23		422	422	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xvtoi_27		422	422	422	vtoi
Xigenebind_6		422	422	422	422	igenebind
Xmm_0		422	422	422	422	422	422	422	422	mm
Xmm_0		422	422	422	422	422	422	422	422	mm
XinputV_95		513	422	vin
XinputV_3		483	166	vin
XinputV_78		475	422	vin
XinputV_35		487	422	vin
XinputV_69		447	422	vin
XinputV_29		510	422	vin
XinputV_55		494	422	vin
XinputV_34		493	422	vin
XinputV_122		513	422	vin
XinputV_123		494	422	vin
XinputV_33		510	413	vin
XinputV_27		434	422	vin
XinputV_51		491	87	vin
XinputV_60		506	422	vin
XinputV_58		512	422	vin
XinputV_108		508	346	vin
XinputV_71		444	422	vin
XinputV_113		474	422	vin
XinputV_103		492	422	vin
XinputV_5		428	422	vin
XinputV_14		494	422	vin
XinputV_111		465	422	vin
XinputV_78		475	422	vin
XinputV_54		494	422	vin
XinputV_114		513	422	vin
XinputV_77		457	422	vin
XinputV_77		457	422	vin
XinputV_44		452	422	vin
XinputV_8		484	422	vin
XinputV_54		494	422	vin
XinputV_72		503	19	vin
XinputV_114		513	422	vin
XinputV_99		513	422	vin
XinputV_109		480	340	vin
XinputV_104		510	422	vin
XinputV_92		513	422	vin
XinputV_42		496	422	vin
XinputV_22		461	422	vin
XinputV_95		513	422	vin
XinputV_123		494	422	vin
XinputV_91		510	422	vin
XinputV_0		465	422	vin
XinputV_2		441	422	vin
XinputV_20		497	422	vin
XinputV_29		510	422	vin
XinputV_123		494	422	vin
XinputV_104		510	422	vin
XinputV_117		499	422	vin
XinputV_86		507	422	vin
XinputV_8		484	422	vin
XinputV_60		506	422	vin
XinputV_95		513	422	vin
XinputV_118		513	422	vin
XinputV_7		484	422	vin
XinputV_114		513	422	vin
XinputV_123		494	422	vin
XinputV_57		485	422	vin
XinputV_122		513	422	vin
XinputV_93		505	422	vin
XinputV_20		497	422	vin
XinputV_8		484	422	vin
XinputV_34		493	422	vin
XinputV_14		494	422	vin
XinputV_102		455	422	vin
XinputV_21		431	327	vin
XinputV_48		450	422	vin
XinputV_118		513	422	vin
XinputV_0		465	422	vin
XinputV_91		510	422	vin
XinputV_64		466	254	vin
XinputV_98		459	62	vin
XinputV_36		506	422	vin
XinputV_76		425	422	vin
XinputV_82		512	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_92		513	422	vin
XinputV_11		463	395	vin
XinputV_6		487	422	vin
XinputV_6		487	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_58		512	422	vin
XinputV_122		513	422	vin
XinputV_99		513	422	vin
XinputV_82		512	422	vin
XinputV_122		513	422	vin
XinputV_122		513	422	vin
XinputV_46		467	422	vin
Xitov_7		422	422	422	itov
Xitov_12		422	422	422	itov
Xitov_16		422	422	422	itov
Xitov_22		422	413	114	itov
Xitov_28		422	422	422	itov
Xitov_24		422	422	422	itov
Xitov_27		422	422	422	itov
Xitov_21		422	422	422	itov
Xitov_5		422	422	422	itov
Xitov_16		422	422	422	itov
Xitov_14		422	422	422	itov
Xitov_21		422	422	422	itov
Xitov_24		422	422	422	itov
Xitov_17		422	422	422	itov
Xitov_25		422	422	422	itov
Xitov_28		422	422	422	itov
Xitov_28		422	422	422	itov
Xitov_17		422	422	422	itov
Xitov_27		422	422	422	itov
Xitov_19		0	422	422	itov
Xitov_28		422	422	422	itov
Xitov_13		422	422	422	itov
Xitov_21		422	422	422	itov
Xitov_28		422	422	422	itov
Xitov_13		422	422	422	itov
Xitov_28		422	422	422	itov
Xitov_27		422	422	422	itov
Xitov_16		422	422	422	itov
Xitov_13		422	422	422	itov
Xitov_5		422	422	422	itov
Xiadd_2		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_12		422	104	11	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_3		422	422	422	422	422	iadd
Xiadd_1		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_0		422	97	422	422	29	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_4		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_28		422	422	422	422	422	iadd
Xiadd_2		422	422	422	422	422	iadd
Xiadd_8		422	422	422	422	422	iadd
Xiadd_28		422	422	422	422	422	iadd
Xiadd_26		422	422	422	422	422	iadd
Xiadd_16		422	387	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_4		422	422	422	422	422	iadd
Xiadd_27		422	422	422	422	422	iadd
Xiadd_20		422	422	422	422	422	iadd
XoutputI_4		422	479	iout
XoutputI_0		422	487	iout
XoutputI_2		422	454	iout
XoutputI_1		29	427	iout
XoutputI_0		422	487	iout
XoutputI_7		422	496	iout
XoutputI_6		422	514	iout
XoutputI_7		422	496	iout
