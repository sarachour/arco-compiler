
*@output LacLp
*@args 141,V
*
*@input TetRp
Iin_TetRp_37		140	0	DC	1.
*
*@input LacLm_0
Vin_LacLm_0_36		140	0	DC	1.
*
*@output TetRp
*@args 139,V
*
*@input TRTetR
Vin_TRTetR_34		139	0	DC	1.
*
*@input clp_0
Vin_clp_0_33		138	0	DC	1.
*
*constant value 752.57498916
Vcst32		137	0	DC	752.57498916
*
*@input TRLacL
Vin_TRLacL_31		136	0	DC	1.
*
*@input clm
Vin_clm_30		135	0	DC	1.
*
*constant value 1.5051499783
Vcst29		135	0	DC	1.5051499783
*
*constant value 0.
Vcst28		135	0	DC	0.
*
*constant value 0.0005
Icst27		134	0	DC	0.0005
*
*@input clp
Iin_clp_26		133	0	DC	1.
*
*@input LacLp
Iin_LacLp_25		132	0	DC	1.
*
*@output LacLm
*@args 131,V
*
*@output TetRm
*@args 130,V
*
*@input KM
Iin_KM_22		129	0	DC	1.
*
*@output TRLacL
*@args 128,I
*
*@output clp
*@args 127,V
*
*constant value 1.
Vcst19		126	0	DC	1.
*
*@input LacLp_0
Vin_LacLp_0_18		125	0	DC	1.
*
*@input TRclp
Vin_TRclp_17		125	0	DC	1.
*
*constant value 0.0332192809489
Vcst16		124	0	DC	0.0332192809489
*
*@input TetRm_0
Vin_TetRm_0_15		123	0	DC	1.
*
*@input TetRm
Vin_TetRm_14		123	0	DC	1.
*
*@input LacLm
Iin_LacLm_13		122	0	DC	1.
*
*@input clm_0
Vin_clm_0_12		122	0	DC	1.
*
*constant value 0.00132877123795
Vcst11		121	0	DC	0.00132877123795
*
*constant value 0.
Icst10		120	0	DC	0.
*
*@output clm
*@args 119,V
*
*constant value 0.4995
Icst8		118	0	DC	0.4995
*
*@output TRclp
*@args 117,I
*
*@output TRTetR
*@args 116,I
*
*constant value 2.
Vcst5		116	0	DC	2.
*
*@input TetRp_0
Vin_TetRp_0_4		115	0	DC	1.
*
*constant value 0.004
Vcst3		114	0	DC	0.004
*
*constant value 250.
Vcst2		113	0	DC	250.
*
*constant value 0.3010299956
Vcst1		112	0	DC	0.3010299956
*
*@input TetRp
Vin_TetRp_0		111	0	DC	1.
*
*
*
* === Connectivity Schem ==== 
Xvgain_24		1	107	23	107	vgain
Xvgain_5		5	107	105	107	vgain
Xvgain_38		107	105	105	107	vgain
Xvgain_38		107	105	105	107	vgain
Xvgain_1		5	107	106	69	vgain
XinputI_3		133	36	iin
XinputI_22		140	38	iin
XinputI_8		134	31	iin
XinputI_11		120	12	iin
XinputI_7		118	90	iin
XinputI_2		132	59	iin
XinputI_19		129	16	iin
XinputI_0		122	49	iin
XoutputV_1		24	127	vout
XoutputV_38		105	131	vout
XoutputV_7		17	130	vout
XoutputV_29		105	139	vout
XoutputV_27		19	141	vout
XoutputV_46		61	119	vout
Xvadd_3		107	107	107	81	0	24	109	vadd
Xvadd_0		107	107	107	105	0	105	105	vadd
Xvadd_30		107	107	107	105	0	17	91	vadd
Xvadd_0		107	107	107	105	0	105	105	vadd
Xvadd_14		75	107	107	81	0	19	53	vadd
Xvadd_21		107	69	107	23	0	61	105	vadd
Xihill_0		90	36	105	16	0	57	ihill
Xihill_1		90	38	105	16	0	34	ihill
Xihill_4		90	59	105	16	0	40	ihill
XinputV_2		137	1	vin
XinputV_41		135	23	vin
XinputV_39		138	109	vin
XinputV_11		140	105	vin
XinputV_33		113	5	vin
XinputV_11		140	105	vin
XinputV_55		135	105	vin
XinputV_73		139	105	vin
XinputV_72		135	107	vin
XinputV_73		139	105	vin
XinputV_69		123	91	vin
XinputV_27		114	105	vin
XinputV_73		139	105	vin
XinputV_72		135	107	vin
XinputV_73		139	105	vin
XinputV_5		111	105	vin
XinputV_55		135	105	vin
XinputV_34		112	81	vin
XinputV_67		125	53	vin
XinputV_46		125	106	vin
XinputV_73		139	105	vin
XinputV_46		125	106	vin
Xitov_11		49	106	75	itov
Xiadd_5		31	57	12	12	63	iadd
Xiadd_17		31	34	12	12	47	iadd
Xiadd_10		31	40	12	12	73	iadd
XoutputI_0		63	117	iout
XoutputI_7		47	116	iout
XoutputI_6		73	128	iout
